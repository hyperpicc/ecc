//Multiplication level4
//April 21, 2009
//Yu Zhang
//yu.zhang100@gmail.com
//verified: y
module level4(L4_A, L4_B, L4_C);
			input 	[177:0]L4_A;
			input 	[177:0]L4_B;
			output 	[193:0]L4_C;
			
			
			assign L4_C[0] = L4_A[0];
			assign L4_C[1] = L4_A[1];
			assign L4_C[2] = L4_A[2];
			assign L4_C[3] = L4_A[3];
			assign L4_C[4] = L4_A[4];
			assign L4_C[5] = L4_A[5];
			assign L4_C[6] = L4_A[6];
			assign L4_C[7] = L4_A[7];
			assign L4_C[8] = L4_A[8];
			assign L4_C[9] = L4_A[9];
			assign L4_C[10] = L4_A[10];
			assign L4_C[11] = L4_A[11];
			assign L4_C[12] = L4_A[12];
			assign L4_C[13] = L4_A[13];
			assign L4_C[14] = L4_A[14];
			assign L4_C[15] = L4_A[15];
			assign L4_C[16] = L4_A[16] ^ L4_B[0];
			assign L4_C[17] = L4_A[17] ^ L4_B[1];
			assign L4_C[18] = L4_A[18] ^ L4_B[2];
			assign L4_C[19] = L4_A[19] ^ L4_B[3];
			assign L4_C[20] = L4_A[20] ^ L4_B[4];
			assign L4_C[21] = L4_A[21] ^ L4_B[5];
			assign L4_C[22] = L4_A[22] ^ L4_B[6];
			assign L4_C[23] = L4_A[23] ^ L4_B[7];
			assign L4_C[24] = L4_A[24] ^ L4_B[8];
			assign L4_C[25] = L4_A[25] ^ L4_B[9];
			assign L4_C[26] = L4_A[26] ^ L4_B[10];
			assign L4_C[27] = L4_A[27] ^ L4_B[11];
			assign L4_C[28] = L4_A[28] ^ L4_B[12];
			assign L4_C[29] = L4_A[29] ^ L4_B[13];
			assign L4_C[30] = L4_A[30] ^ L4_B[14];
			assign L4_C[31] = L4_A[31] ^ L4_B[15];
			assign L4_C[32] = L4_A[32] ^ L4_B[16];
			assign L4_C[33] = L4_A[33] ^ L4_B[17];
			assign L4_C[34] = L4_A[34] ^ L4_B[18];
			assign L4_C[35] = L4_A[35] ^ L4_B[19];
			assign L4_C[36] = L4_A[36] ^ L4_B[20];
			assign L4_C[37] = L4_A[37] ^ L4_B[21];
			assign L4_C[38] = L4_A[38] ^ L4_B[22];
			assign L4_C[39] = L4_A[39] ^ L4_B[23];
			assign L4_C[40] = L4_A[40] ^ L4_B[24];
			assign L4_C[41] = L4_A[41] ^ L4_B[25];
			assign L4_C[42] = L4_A[42] ^ L4_B[26];
			assign L4_C[43] = L4_A[43] ^ L4_B[27];
			assign L4_C[44] = L4_A[44] ^ L4_B[28];
			assign L4_C[45] = L4_A[45] ^ L4_B[29];
			assign L4_C[46] = L4_A[46] ^ L4_B[30];
			assign L4_C[47] = L4_A[47] ^ L4_B[31];
			assign L4_C[48] = L4_A[48] ^ L4_B[32];
			assign L4_C[49] = L4_A[49] ^ L4_B[33];
			assign L4_C[50] = L4_A[50] ^ L4_B[34];
			assign L4_C[51] = L4_A[51] ^ L4_B[35];
			assign L4_C[52] = L4_A[52] ^ L4_B[36];
			assign L4_C[53] = L4_A[53] ^ L4_B[37];
			assign L4_C[54] = L4_A[54] ^ L4_B[38];
			assign L4_C[55] = L4_A[55] ^ L4_B[39];
			assign L4_C[56] = L4_A[56] ^ L4_B[40];
			assign L4_C[57] = L4_A[57] ^ L4_B[41];
			assign L4_C[58] = L4_A[58] ^ L4_B[42];
			assign L4_C[59] = L4_A[59] ^ L4_B[43];
			assign L4_C[60] = L4_A[60] ^ L4_B[44];
			assign L4_C[61] = L4_A[61] ^ L4_B[45];
			assign L4_C[62] = L4_A[62] ^ L4_B[46];
			assign L4_C[63] = L4_A[63] ^ L4_B[47];
			assign L4_C[64] = L4_A[64] ^ L4_B[48];
			assign L4_C[65] = L4_A[65] ^ L4_B[49];
			assign L4_C[66] = L4_A[66] ^ L4_B[50];
			assign L4_C[67] = L4_A[67] ^ L4_B[51];
			assign L4_C[68] = L4_A[68] ^ L4_B[52];
			assign L4_C[69] = L4_A[69] ^ L4_B[53];
			assign L4_C[70] = L4_A[70] ^ L4_B[54];
			assign L4_C[71] = L4_A[71] ^ L4_B[55];
			assign L4_C[72] = L4_A[72] ^ L4_B[56];
			assign L4_C[73] = L4_A[73] ^ L4_B[57];
			assign L4_C[74] = L4_A[74] ^ L4_B[58];
			assign L4_C[75] = L4_A[75] ^ L4_B[59];
			assign L4_C[76] = L4_A[76] ^ L4_B[60];
			assign L4_C[77] = L4_A[77] ^ L4_B[61];
			assign L4_C[78] = L4_A[78] ^ L4_B[62];
			assign L4_C[79] = L4_A[79] ^ L4_B[63];
			assign L4_C[80] = L4_A[80] ^ L4_B[64];
			assign L4_C[81] = L4_A[81] ^ L4_B[65];
			assign L4_C[82] = L4_A[82] ^ L4_B[66];
			assign L4_C[83] = L4_A[83] ^ L4_B[67];
			assign L4_C[84] = L4_A[84] ^ L4_B[68];
			assign L4_C[85] = L4_A[85] ^ L4_B[69];
			assign L4_C[86] = L4_A[86] ^ L4_B[70];
			assign L4_C[87] = L4_A[87] ^ L4_B[71];
			assign L4_C[88] = L4_A[88] ^ L4_B[72];
			assign L4_C[89] = L4_A[89] ^ L4_B[73];
			assign L4_C[90] = L4_A[90] ^ L4_B[74];
			assign L4_C[91] = L4_A[91] ^ L4_B[75];
			assign L4_C[92] = L4_A[92] ^ L4_B[76];
			assign L4_C[93] = L4_A[93] ^ L4_B[77];
			assign L4_C[94] = L4_A[94] ^ L4_B[78];
			assign L4_C[95] = L4_A[95] ^ L4_B[79];
			assign L4_C[96] = L4_A[96] ^ L4_B[80];
			assign L4_C[97] = L4_A[97] ^ L4_B[81];
			assign L4_C[98] = L4_A[98] ^ L4_B[82];
			assign L4_C[99] = L4_A[99] ^ L4_B[83];
			assign L4_C[100] = L4_A[100] ^ L4_B[84];
			assign L4_C[101] = L4_A[101] ^ L4_B[85];
			assign L4_C[102] = L4_A[102] ^ L4_B[86];
			assign L4_C[103] = L4_A[103] ^ L4_B[87];
			assign L4_C[104] = L4_A[104] ^ L4_B[88];
			assign L4_C[105] = L4_A[105] ^ L4_B[89];
			assign L4_C[106] = L4_A[106] ^ L4_B[90];
			assign L4_C[107] = L4_A[107] ^ L4_B[91];
			assign L4_C[108] = L4_A[108] ^ L4_B[92];
			assign L4_C[109] = L4_A[109] ^ L4_B[93];
			assign L4_C[110] = L4_A[110] ^ L4_B[94];
			assign L4_C[111] = L4_A[111] ^ L4_B[95];
			assign L4_C[112] = L4_A[112] ^ L4_B[96];
			assign L4_C[113] = L4_A[113] ^ L4_B[97];
			assign L4_C[114] = L4_A[114] ^ L4_B[98];
			assign L4_C[115] = L4_A[115] ^ L4_B[99];
			assign L4_C[116] = L4_A[116] ^ L4_B[100];
			assign L4_C[117] = L4_A[117] ^ L4_B[101];
			assign L4_C[118] = L4_A[118] ^ L4_B[102];
			assign L4_C[119] = L4_A[119] ^ L4_B[103];
			assign L4_C[120] = L4_A[120] ^ L4_B[104];
			assign L4_C[121] = L4_A[121] ^ L4_B[105];
			assign L4_C[122] = L4_A[122] ^ L4_B[106];
			assign L4_C[123] = L4_A[123] ^ L4_B[107];
			assign L4_C[124] = L4_A[124] ^ L4_B[108];
			assign L4_C[125] = L4_A[125] ^ L4_B[109];
			assign L4_C[126] = L4_A[126] ^ L4_B[110];
			assign L4_C[127] = L4_A[127] ^ L4_B[111];
			assign L4_C[128] = L4_A[128] ^ L4_B[112];
			assign L4_C[129] = L4_A[129] ^ L4_B[113];
			assign L4_C[130] = L4_A[130] ^ L4_B[114];
			assign L4_C[131] = L4_A[131] ^ L4_B[115];
			assign L4_C[132] = L4_A[132] ^ L4_B[116];
			assign L4_C[133] = L4_A[133] ^ L4_B[117];
			assign L4_C[134] = L4_A[134] ^ L4_B[118];
			assign L4_C[135] = L4_A[135] ^ L4_B[119];
			assign L4_C[136] = L4_A[136] ^ L4_B[120];
			assign L4_C[137] = L4_A[137] ^ L4_B[121];
			assign L4_C[138] = L4_A[138] ^ L4_B[122];
			assign L4_C[139] = L4_A[139] ^ L4_B[123];
			assign L4_C[140] = L4_A[140] ^ L4_B[124];
			assign L4_C[141] = L4_A[141] ^ L4_B[125];
			assign L4_C[142] = L4_A[142] ^ L4_B[126];
			assign L4_C[143] = L4_A[143] ^ L4_B[127];
			assign L4_C[144] = L4_A[144] ^ L4_B[128];
			assign L4_C[145] = L4_A[145] ^ L4_B[129];
			assign L4_C[146] = L4_A[146] ^ L4_B[130];
			assign L4_C[147] = L4_A[147] ^ L4_B[131];
			assign L4_C[148] = L4_A[148] ^ L4_B[132];
			assign L4_C[149] = L4_A[149] ^ L4_B[133];
			assign L4_C[150] = L4_A[150] ^ L4_B[134];
			assign L4_C[151] = L4_A[151] ^ L4_B[135];
			assign L4_C[152] = L4_A[152] ^ L4_B[136];
			assign L4_C[153] = L4_A[153] ^ L4_B[137];
			assign L4_C[154] = L4_A[154] ^ L4_B[138];
			assign L4_C[155] = L4_A[155] ^ L4_B[139];
			assign L4_C[156] = L4_A[156] ^ L4_B[140];
			assign L4_C[157] = L4_A[157] ^ L4_B[141];
			assign L4_C[158] = L4_A[158] ^ L4_B[142];
			assign L4_C[159] = L4_A[159] ^ L4_B[143];
			assign L4_C[160] = L4_A[160] ^ L4_B[144];
			assign L4_C[161] = L4_A[161] ^ L4_B[145];
			assign L4_C[162] = L4_A[162] ^ L4_B[146];
			assign L4_C[163] = L4_A[163] ^ L4_B[147];
			assign L4_C[164] = L4_A[164] ^ L4_B[148];
			assign L4_C[165] = L4_A[165] ^ L4_B[149];
			assign L4_C[166] = L4_A[166] ^ L4_B[150];
			assign L4_C[167] = L4_A[167] ^ L4_B[151];
			assign L4_C[168] = L4_A[168] ^ L4_B[152];
			assign L4_C[169] = L4_A[169] ^ L4_B[153];
			assign L4_C[170] = L4_A[170] ^ L4_B[154];
			assign L4_C[171] = L4_A[171] ^ L4_B[155];
			assign L4_C[172] = L4_A[172] ^ L4_B[156];
			assign L4_C[173] = L4_A[173] ^ L4_B[157];
			assign L4_C[174] = L4_A[174] ^ L4_B[158];
			assign L4_C[175] = L4_A[175] ^ L4_B[159];
			assign L4_C[176] = L4_A[176] ^ L4_B[160];
			assign L4_C[177] = L4_A[177] ^ L4_B[161];		
			assign L4_C[178] = L4_B[162];
			assign L4_C[179] = L4_B[163];
			assign L4_C[180] = L4_B[164];
			assign L4_C[181] = L4_B[165];
			assign L4_C[182] = L4_B[166];
			assign L4_C[183] = L4_B[167];
			assign L4_C[184] = L4_B[168];
			assign L4_C[185] = L4_B[169];
			assign L4_C[186] = L4_B[170];
			assign L4_C[187] = L4_B[171];
			assign L4_C[188] = L4_B[172];
			assign L4_C[189] = L4_B[173];
			assign L4_C[190] = L4_B[174];
			assign L4_C[191] = L4_B[175];
			assign L4_C[192] = L4_B[176];
			assign L4_C[193] = L4_B[177];
endmodule
