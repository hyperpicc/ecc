//Multiplication level2
//April 21, 2009
//Yu Zhang
//yu.zhang100@gmail.com
//verified: y
module level2(L2_A, L2_B, L2_C);
			input 	[165:0]L2_A;
			input 	[165:0]L2_B;
			output 	[169:0]L2_C;
				
				
				assign L2_C[0] = L2_A[0] ;
				assign L2_C[1] = L2_A[1] ;
				assign L2_C[2] = L2_A[2] ;
				assign L2_C[3] = L2_A[3] ;
			  assign L2_C[4] = L2_A[4] ^ L2_B[0];
				assign L2_C[5] = L2_A[5] ^ L2_B[1];
				assign L2_C[6] = L2_A[6] ^ L2_B[2];
				assign L2_C[7] = L2_A[7] ^ L2_B[3];
				assign L2_C[8] = L2_A[8] ^ L2_B[4];
				assign L2_C[9] = L2_A[9] ^ L2_B[5];
				assign L2_C[10] = L2_A[10] ^ L2_B[6];
				assign L2_C[11] = L2_A[11] ^ L2_B[7];
				assign L2_C[12] = L2_A[12] ^ L2_B[8];
				assign L2_C[13] = L2_A[13] ^ L2_B[9];
				assign L2_C[14] = L2_A[14] ^ L2_B[10];
				assign L2_C[15] = L2_A[15] ^ L2_B[11];
				assign L2_C[16] = L2_A[16] ^ L2_B[12];
				assign L2_C[17] = L2_A[17] ^ L2_B[13];
				assign L2_C[18] = L2_A[18] ^ L2_B[14];
				assign L2_C[19] = L2_A[19] ^ L2_B[15];
				assign L2_C[20] = L2_A[20] ^ L2_B[16];
				assign L2_C[21] = L2_A[21] ^ L2_B[17];
				assign L2_C[22] = L2_A[22] ^ L2_B[18];
				assign L2_C[23] = L2_A[23] ^ L2_B[19];
				assign L2_C[24] = L2_A[24] ^ L2_B[20];
				assign L2_C[25] = L2_A[25] ^ L2_B[21];
				assign L2_C[26] = L2_A[26] ^ L2_B[22];
				assign L2_C[27] = L2_A[27] ^ L2_B[23];
				assign L2_C[28] = L2_A[28] ^ L2_B[24];
				assign L2_C[29] = L2_A[29] ^ L2_B[25];
				assign L2_C[30] = L2_A[30] ^ L2_B[26];
				assign L2_C[31] = L2_A[31] ^ L2_B[27];
				assign L2_C[32] = L2_A[32] ^ L2_B[28];
				assign L2_C[33] = L2_A[33] ^ L2_B[29];
				assign L2_C[34] = L2_A[34] ^ L2_B[30];
				assign L2_C[35] = L2_A[35] ^ L2_B[31];
				assign L2_C[36] = L2_A[36] ^ L2_B[32];
				assign L2_C[37] = L2_A[37] ^ L2_B[33];
				assign L2_C[38] = L2_A[38] ^ L2_B[34];
				assign L2_C[39] = L2_A[39] ^ L2_B[35];
				assign L2_C[40] = L2_A[40] ^ L2_B[36];
				assign L2_C[41] = L2_A[41] ^ L2_B[37];
				assign L2_C[42] = L2_A[42] ^ L2_B[38];
				assign L2_C[43] = L2_A[43] ^ L2_B[39];
				assign L2_C[44] = L2_A[44] ^ L2_B[40];
				assign L2_C[45] = L2_A[45] ^ L2_B[41];
				assign L2_C[46] = L2_A[46] ^ L2_B[42];
				assign L2_C[47] = L2_A[47] ^ L2_B[43];
				assign L2_C[48] = L2_A[48] ^ L2_B[44];
				assign L2_C[49] = L2_A[49] ^ L2_B[45];
				assign L2_C[50] = L2_A[50] ^ L2_B[46];
				assign L2_C[51] = L2_A[51] ^ L2_B[47];
				assign L2_C[52] = L2_A[52] ^ L2_B[48];
				assign L2_C[53] = L2_A[53] ^ L2_B[49];
				assign L2_C[54] = L2_A[54] ^ L2_B[50];
				assign L2_C[55] = L2_A[55] ^ L2_B[51];
				assign L2_C[56] = L2_A[56] ^ L2_B[52];
				assign L2_C[57] = L2_A[57] ^ L2_B[53];
				assign L2_C[58] = L2_A[58] ^ L2_B[54];
				assign L2_C[59] = L2_A[59] ^ L2_B[55];
				assign L2_C[60] = L2_A[60] ^ L2_B[56];
				assign L2_C[61] = L2_A[61] ^ L2_B[57];
				assign L2_C[62] = L2_A[62] ^ L2_B[58];
				assign L2_C[63] = L2_A[63] ^ L2_B[59];
				assign L2_C[64] = L2_A[64] ^ L2_B[60];
				assign L2_C[65] = L2_A[65] ^ L2_B[61];
				assign L2_C[66] = L2_A[66] ^ L2_B[62];
				assign L2_C[67] = L2_A[67] ^ L2_B[63];
				assign L2_C[68] = L2_A[68] ^ L2_B[64];
				assign L2_C[69] = L2_A[69] ^ L2_B[65];
				assign L2_C[70] = L2_A[70] ^ L2_B[66];
				assign L2_C[71] = L2_A[71] ^ L2_B[67];
				assign L2_C[72] = L2_A[72] ^ L2_B[68];
				assign L2_C[73] = L2_A[73] ^ L2_B[69];
				assign L2_C[74] = L2_A[74] ^ L2_B[70];
				assign L2_C[75] = L2_A[75] ^ L2_B[71];
				assign L2_C[76] = L2_A[76] ^ L2_B[72];
				assign L2_C[77] = L2_A[77] ^ L2_B[73];
				assign L2_C[78] = L2_A[78] ^ L2_B[74];
				assign L2_C[79] = L2_A[79] ^ L2_B[75];
				assign L2_C[80] = L2_A[80] ^ L2_B[76];
				assign L2_C[81] = L2_A[81] ^ L2_B[77];
				assign L2_C[82] = L2_A[82] ^ L2_B[78];
				assign L2_C[83] = L2_A[83] ^ L2_B[79];
				assign L2_C[84] = L2_A[84] ^ L2_B[80];
				assign L2_C[85] = L2_A[85] ^ L2_B[81];
				assign L2_C[86] = L2_A[86] ^ L2_B[82];
				assign L2_C[87] = L2_A[87] ^ L2_B[83];
				assign L2_C[88] = L2_A[88] ^ L2_B[84];
				assign L2_C[89] = L2_A[89] ^ L2_B[85];
				assign L2_C[90] = L2_A[90] ^ L2_B[86];
				assign L2_C[91] = L2_A[91] ^ L2_B[87];
				assign L2_C[92] = L2_A[92] ^ L2_B[88];
				assign L2_C[93] = L2_A[93] ^ L2_B[89];
				assign L2_C[94] = L2_A[94] ^ L2_B[90];
				assign L2_C[95] = L2_A[95] ^ L2_B[91];
				assign L2_C[96] = L2_A[96] ^ L2_B[92];
				assign L2_C[97] = L2_A[97] ^ L2_B[93];
				assign L2_C[98] = L2_A[98] ^ L2_B[94];
				assign L2_C[99] = L2_A[99] ^ L2_B[95];
				assign L2_C[100] = L2_A[100] ^ L2_B[96];
				assign L2_C[101] = L2_A[101] ^ L2_B[97];
				assign L2_C[102] = L2_A[102] ^ L2_B[98];
				assign L2_C[103] = L2_A[103] ^ L2_B[99];
				assign L2_C[104] = L2_A[104] ^ L2_B[100];
				assign L2_C[105] = L2_A[105] ^ L2_B[101];
				assign L2_C[106] = L2_A[106] ^ L2_B[102];
				assign L2_C[107] = L2_A[107] ^ L2_B[103];
				assign L2_C[108] = L2_A[108] ^ L2_B[104];
				assign L2_C[109] = L2_A[109] ^ L2_B[105];
				assign L2_C[110] = L2_A[110] ^ L2_B[106];
				assign L2_C[111] = L2_A[111] ^ L2_B[107];
				assign L2_C[112] = L2_A[112] ^ L2_B[108];
				assign L2_C[113] = L2_A[113] ^ L2_B[109];
				assign L2_C[114] = L2_A[114] ^ L2_B[110];
				assign L2_C[115] = L2_A[115] ^ L2_B[111];
				assign L2_C[116] = L2_A[116] ^ L2_B[112];
				assign L2_C[117] = L2_A[117] ^ L2_B[113];
				assign L2_C[118] = L2_A[118] ^ L2_B[114];
				assign L2_C[119] = L2_A[119] ^ L2_B[115];
				assign L2_C[120] = L2_A[120] ^ L2_B[116];
				assign L2_C[121] = L2_A[121] ^ L2_B[117];
				assign L2_C[122] = L2_A[122] ^ L2_B[118];
				assign L2_C[123] = L2_A[123] ^ L2_B[119];
				assign L2_C[124] = L2_A[124] ^ L2_B[120];
				assign L2_C[125] = L2_A[125] ^ L2_B[121];
				assign L2_C[126] = L2_A[126] ^ L2_B[122];
				assign L2_C[127] = L2_A[127] ^ L2_B[123];
				assign L2_C[128] = L2_A[128] ^ L2_B[124];
				assign L2_C[129] = L2_A[129] ^ L2_B[125];
				assign L2_C[130] = L2_A[130] ^ L2_B[126];
				assign L2_C[131] = L2_A[131] ^ L2_B[127];
				assign L2_C[132] = L2_A[132] ^ L2_B[128];
				assign L2_C[133] = L2_A[133] ^ L2_B[129];
				assign L2_C[134] = L2_A[134] ^ L2_B[130];
				assign L2_C[135] = L2_A[135] ^ L2_B[131];
				assign L2_C[136] = L2_A[136] ^ L2_B[132];
				assign L2_C[137] = L2_A[137] ^ L2_B[133];
				assign L2_C[138] = L2_A[138] ^ L2_B[134];
				assign L2_C[139] = L2_A[139] ^ L2_B[135];
				assign L2_C[140] = L2_A[140] ^ L2_B[136];
				assign L2_C[141] = L2_A[141] ^ L2_B[137];
				assign L2_C[142] = L2_A[142] ^ L2_B[138];
				assign L2_C[143] = L2_A[143] ^ L2_B[139];
				assign L2_C[144] = L2_A[144] ^ L2_B[140];
				assign L2_C[145] = L2_A[145] ^ L2_B[141];
				assign L2_C[146] = L2_A[146] ^ L2_B[142];
				assign L2_C[147] = L2_A[147] ^ L2_B[143];
				assign L2_C[148] = L2_A[148] ^ L2_B[144];
				assign L2_C[149] = L2_A[149] ^ L2_B[145];
				assign L2_C[150] = L2_A[150] ^ L2_B[146];
				assign L2_C[151] = L2_A[151] ^ L2_B[147];
				assign L2_C[152] = L2_A[152] ^ L2_B[148];
				assign L2_C[153] = L2_A[153] ^ L2_B[149];
				assign L2_C[154] = L2_A[154] ^ L2_B[150];
				assign L2_C[155] = L2_A[155] ^ L2_B[151];
				assign L2_C[156] = L2_A[156] ^ L2_B[152];
				assign L2_C[157] = L2_A[157] ^ L2_B[153];
				assign L2_C[158] = L2_A[158] ^ L2_B[154];
				assign L2_C[159] = L2_A[159] ^ L2_B[155];
				assign L2_C[160] = L2_A[160] ^ L2_B[156];
				assign L2_C[161] = L2_A[161] ^ L2_B[157];
				assign L2_C[162] = L2_A[162] ^ L2_B[158];
				assign L2_C[163] = L2_A[163] ^ L2_B[159];
				assign L2_C[164] = L2_A[164] ^ L2_B[160];
				assign L2_C[165] = L2_A[165] ^ L2_B[161];
				assign L2_C[166] = L2_B[162];
				assign L2_C[167] = L2_B[163];
				assign L2_C[168] = L2_B[164];
				assign L2_C[169] = L2_B[165];			
				
			endmodule
