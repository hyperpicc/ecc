//Multiplication level0
//April 21, 2009
//Yu Zhang
//yu.zhang100@gmail.com
//verified: y
			module level0(L0_A, L0_B, L0_C);
			input 	[1:0]L0_A;
			input 	[162:0]L0_B;
			output 	[163:0]L0_C;


			
			assign L0_C[0] = L0_A[0] & L0_B[0];
			assign L0_C[1] = L0_A[0] & L0_B[1] ^ L0_A[1] & L0_B[0];
			assign L0_C[2] = L0_A[0] & L0_B[2] ^ L0_A[1] & L0_B[1];
			assign L0_C[3] = L0_A[0] & L0_B[3] ^ L0_A[1] & L0_B[2];
			assign L0_C[4] = L0_A[0] & L0_B[4] ^ L0_A[1] & L0_B[3];
			assign L0_C[5] = L0_A[0] & L0_B[5] ^ L0_A[1] & L0_B[4];
			assign L0_C[6] = L0_A[0] & L0_B[6] ^ L0_A[1] & L0_B[5];
			assign L0_C[7] = L0_A[0] & L0_B[7] ^ L0_A[1] & L0_B[6];
			assign L0_C[8] = L0_A[0] & L0_B[8] ^ L0_A[1] & L0_B[7];
			assign L0_C[9] = L0_A[0] & L0_B[9] ^ L0_A[1] & L0_B[8];
			assign L0_C[10] = L0_A[0] & L0_B[10] ^ L0_A[1] & L0_B[9];
			assign L0_C[11] = L0_A[0] & L0_B[11] ^ L0_A[1] & L0_B[10];
			assign L0_C[12] = L0_A[0] & L0_B[12] ^ L0_A[1] & L0_B[11];
			assign L0_C[13] = L0_A[0] & L0_B[13] ^ L0_A[1] & L0_B[12];
			assign L0_C[14] = L0_A[0] & L0_B[14] ^ L0_A[1] & L0_B[13];
			assign L0_C[15] = L0_A[0] & L0_B[15] ^ L0_A[1] & L0_B[14];
			assign L0_C[16] = L0_A[0] & L0_B[16] ^ L0_A[1] & L0_B[15];
			assign L0_C[17] = L0_A[0] & L0_B[17] ^ L0_A[1] & L0_B[16];
			assign L0_C[18] = L0_A[0] & L0_B[18] ^ L0_A[1] & L0_B[17];
			assign L0_C[19] = L0_A[0] & L0_B[19] ^ L0_A[1] & L0_B[18];
			assign L0_C[20] = L0_A[0] & L0_B[20] ^ L0_A[1] & L0_B[19];
			assign L0_C[21] = L0_A[0] & L0_B[21] ^ L0_A[1] & L0_B[20];
			assign L0_C[22] = L0_A[0] & L0_B[22] ^ L0_A[1] & L0_B[21];
			assign L0_C[23] = L0_A[0] & L0_B[23] ^ L0_A[1] & L0_B[22];
			assign L0_C[24] = L0_A[0] & L0_B[24] ^ L0_A[1] & L0_B[23];
			assign L0_C[25] = L0_A[0] & L0_B[25] ^ L0_A[1] & L0_B[24];
			assign L0_C[26] = L0_A[0] & L0_B[26] ^ L0_A[1] & L0_B[25];
			assign L0_C[27] = L0_A[0] & L0_B[27] ^ L0_A[1] & L0_B[26];
			assign L0_C[28] = L0_A[0] & L0_B[28] ^ L0_A[1] & L0_B[27];
			assign L0_C[29] = L0_A[0] & L0_B[29] ^ L0_A[1] & L0_B[28];
			assign L0_C[30] = L0_A[0] & L0_B[30] ^ L0_A[1] & L0_B[29];
			assign L0_C[31] = L0_A[0] & L0_B[31] ^ L0_A[1] & L0_B[30];
			assign L0_C[32] = L0_A[0] & L0_B[32] ^ L0_A[1] & L0_B[31];
			assign L0_C[33] = L0_A[0] & L0_B[33] ^ L0_A[1] & L0_B[32];
			assign L0_C[34] = L0_A[0] & L0_B[34] ^ L0_A[1] & L0_B[33];
			assign L0_C[35] = L0_A[0] & L0_B[35] ^ L0_A[1] & L0_B[34];
			assign L0_C[36] = L0_A[0] & L0_B[36] ^ L0_A[1] & L0_B[35];
			assign L0_C[37] = L0_A[0] & L0_B[37] ^ L0_A[1] & L0_B[36];
			assign L0_C[38] = L0_A[0] & L0_B[38] ^ L0_A[1] & L0_B[37];
			assign L0_C[39] = L0_A[0] & L0_B[39] ^ L0_A[1] & L0_B[38];
			assign L0_C[40] = L0_A[0] & L0_B[40] ^ L0_A[1] & L0_B[39];
			assign L0_C[41] = L0_A[0] & L0_B[41] ^ L0_A[1] & L0_B[40];
			assign L0_C[42] = L0_A[0] & L0_B[42] ^ L0_A[1] & L0_B[41];
			assign L0_C[43] = L0_A[0] & L0_B[43] ^ L0_A[1] & L0_B[42];
			assign L0_C[44] = L0_A[0] & L0_B[44] ^ L0_A[1] & L0_B[43];
			assign L0_C[45] = L0_A[0] & L0_B[45] ^ L0_A[1] & L0_B[44];
			assign L0_C[46] = L0_A[0] & L0_B[46] ^ L0_A[1] & L0_B[45];
			assign L0_C[47] = L0_A[0] & L0_B[47] ^ L0_A[1] & L0_B[46];
			assign L0_C[48] = L0_A[0] & L0_B[48] ^ L0_A[1] & L0_B[47];
			assign L0_C[49] = L0_A[0] & L0_B[49] ^ L0_A[1] & L0_B[48];
			assign L0_C[50] = L0_A[0] & L0_B[50] ^ L0_A[1] & L0_B[49];
			assign L0_C[51] = L0_A[0] & L0_B[51] ^ L0_A[1] & L0_B[50];
			assign L0_C[52] = L0_A[0] & L0_B[52] ^ L0_A[1] & L0_B[51];
			assign L0_C[53] = L0_A[0] & L0_B[53] ^ L0_A[1] & L0_B[52];
			assign L0_C[54] = L0_A[0] & L0_B[54] ^ L0_A[1] & L0_B[53];
			assign L0_C[55] = L0_A[0] & L0_B[55] ^ L0_A[1] & L0_B[54];
			assign L0_C[56] = L0_A[0] & L0_B[56] ^ L0_A[1] & L0_B[55];
			assign L0_C[57] = L0_A[0] & L0_B[57] ^ L0_A[1] & L0_B[56];
			assign L0_C[58] = L0_A[0] & L0_B[58] ^ L0_A[1] & L0_B[57];
			assign L0_C[59] = L0_A[0] & L0_B[59] ^ L0_A[1] & L0_B[58];
			assign L0_C[60] = L0_A[0] & L0_B[60] ^ L0_A[1] & L0_B[59];
			assign L0_C[61] = L0_A[0] & L0_B[61] ^ L0_A[1] & L0_B[60];
			assign L0_C[62] = L0_A[0] & L0_B[62] ^ L0_A[1] & L0_B[61];
			assign L0_C[63] = L0_A[0] & L0_B[63] ^ L0_A[1] & L0_B[62];
			assign L0_C[64] = L0_A[0] & L0_B[64] ^ L0_A[1] & L0_B[63];
			assign L0_C[65] = L0_A[0] & L0_B[65] ^ L0_A[1] & L0_B[64];
			assign L0_C[66] = L0_A[0] & L0_B[66] ^ L0_A[1] & L0_B[65];
			assign L0_C[67] = L0_A[0] & L0_B[67] ^ L0_A[1] & L0_B[66];
			assign L0_C[68] = L0_A[0] & L0_B[68] ^ L0_A[1] & L0_B[67];
			assign L0_C[69] = L0_A[0] & L0_B[69] ^ L0_A[1] & L0_B[68];
			assign L0_C[70] = L0_A[0] & L0_B[70] ^ L0_A[1] & L0_B[69];
			assign L0_C[71] = L0_A[0] & L0_B[71] ^ L0_A[1] & L0_B[70];
			assign L0_C[72] = L0_A[0] & L0_B[72] ^ L0_A[1] & L0_B[71];
			assign L0_C[73] = L0_A[0] & L0_B[73] ^ L0_A[1] & L0_B[72];
			assign L0_C[74] = L0_A[0] & L0_B[74] ^ L0_A[1] & L0_B[73];
			assign L0_C[75] = L0_A[0] & L0_B[75] ^ L0_A[1] & L0_B[74];
			assign L0_C[76] = L0_A[0] & L0_B[76] ^ L0_A[1] & L0_B[75];
			assign L0_C[77] = L0_A[0] & L0_B[77] ^ L0_A[1] & L0_B[76];
			assign L0_C[78] = L0_A[0] & L0_B[78] ^ L0_A[1] & L0_B[77];
			assign L0_C[79] = L0_A[0] & L0_B[79] ^ L0_A[1] & L0_B[78];
			assign L0_C[80] = L0_A[0] & L0_B[80] ^ L0_A[1] & L0_B[79];
			assign L0_C[81] = L0_A[0] & L0_B[81] ^ L0_A[1] & L0_B[80];
			assign L0_C[82] = L0_A[0] & L0_B[82] ^ L0_A[1] & L0_B[81];
			assign L0_C[83] = L0_A[0] & L0_B[83] ^ L0_A[1] & L0_B[82];
			assign L0_C[84] = L0_A[0] & L0_B[84] ^ L0_A[1] & L0_B[83];
			assign L0_C[85] = L0_A[0] & L0_B[85] ^ L0_A[1] & L0_B[84];
			assign L0_C[86] = L0_A[0] & L0_B[86] ^ L0_A[1] & L0_B[85];
			assign L0_C[87] = L0_A[0] & L0_B[87] ^ L0_A[1] & L0_B[86];
			assign L0_C[88] = L0_A[0] & L0_B[88] ^ L0_A[1] & L0_B[87];
			assign L0_C[89] = L0_A[0] & L0_B[89] ^ L0_A[1] & L0_B[88];
			assign L0_C[90] = L0_A[0] & L0_B[90] ^ L0_A[1] & L0_B[89];
			assign L0_C[91] = L0_A[0] & L0_B[91] ^ L0_A[1] & L0_B[90];
			assign L0_C[92] = L0_A[0] & L0_B[92] ^ L0_A[1] & L0_B[91];
			assign L0_C[93] = L0_A[0] & L0_B[93] ^ L0_A[1] & L0_B[92];
			assign L0_C[94] = L0_A[0] & L0_B[94] ^ L0_A[1] & L0_B[93];
			assign L0_C[95] = L0_A[0] & L0_B[95] ^ L0_A[1] & L0_B[94];
			assign L0_C[96] = L0_A[0] & L0_B[96] ^ L0_A[1] & L0_B[95];
			assign L0_C[97] = L0_A[0] & L0_B[97] ^ L0_A[1] & L0_B[96];
			assign L0_C[98] = L0_A[0] & L0_B[98] ^ L0_A[1] & L0_B[97];
			assign L0_C[99] = L0_A[0] & L0_B[99] ^ L0_A[1] & L0_B[98];
			assign L0_C[100] = L0_A[0] & L0_B[100] ^ L0_A[1] & L0_B[99];
			assign L0_C[101] = L0_A[0] & L0_B[101] ^ L0_A[1] & L0_B[100];
			assign L0_C[102] = L0_A[0] & L0_B[102] ^ L0_A[1] & L0_B[101];
			assign L0_C[103] = L0_A[0] & L0_B[103] ^ L0_A[1] & L0_B[102];
			assign L0_C[104] = L0_A[0] & L0_B[104] ^ L0_A[1] & L0_B[103];
			assign L0_C[105] = L0_A[0] & L0_B[105] ^ L0_A[1] & L0_B[104];
			assign L0_C[106] = L0_A[0] & L0_B[106] ^ L0_A[1] & L0_B[105];
			assign L0_C[107] = L0_A[0] & L0_B[107] ^ L0_A[1] & L0_B[106];
			assign L0_C[108] = L0_A[0] & L0_B[108] ^ L0_A[1] & L0_B[107];
			assign L0_C[109] = L0_A[0] & L0_B[109] ^ L0_A[1] & L0_B[108];
			assign L0_C[110] = L0_A[0] & L0_B[110] ^ L0_A[1] & L0_B[109];
			assign L0_C[111] = L0_A[0] & L0_B[111] ^ L0_A[1] & L0_B[110];
			assign L0_C[112] = L0_A[0] & L0_B[112] ^ L0_A[1] & L0_B[111];
			assign L0_C[113] = L0_A[0] & L0_B[113] ^ L0_A[1] & L0_B[112];
			assign L0_C[114] = L0_A[0] & L0_B[114] ^ L0_A[1] & L0_B[113];
			assign L0_C[115] = L0_A[0] & L0_B[115] ^ L0_A[1] & L0_B[114];
			assign L0_C[116] = L0_A[0] & L0_B[116] ^ L0_A[1] & L0_B[115];
			assign L0_C[117] = L0_A[0] & L0_B[117] ^ L0_A[1] & L0_B[116];
			assign L0_C[118] = L0_A[0] & L0_B[118] ^ L0_A[1] & L0_B[117];
			assign L0_C[119] = L0_A[0] & L0_B[119] ^ L0_A[1] & L0_B[118];
			assign L0_C[120] = L0_A[0] & L0_B[120] ^ L0_A[1] & L0_B[119];
			assign L0_C[121] = L0_A[0] & L0_B[121] ^ L0_A[1] & L0_B[120];
			assign L0_C[122] = L0_A[0] & L0_B[122] ^ L0_A[1] & L0_B[121];
			assign L0_C[123] = L0_A[0] & L0_B[123] ^ L0_A[1] & L0_B[122];
			assign L0_C[124] = L0_A[0] & L0_B[124] ^ L0_A[1] & L0_B[123];
			assign L0_C[125] = L0_A[0] & L0_B[125] ^ L0_A[1] & L0_B[124];
			assign L0_C[126] = L0_A[0] & L0_B[126] ^ L0_A[1] & L0_B[125];
			assign L0_C[127] = L0_A[0] & L0_B[127] ^ L0_A[1] & L0_B[126];
			assign L0_C[128] = L0_A[0] & L0_B[128] ^ L0_A[1] & L0_B[127];
			assign L0_C[129] = L0_A[0] & L0_B[129] ^ L0_A[1] & L0_B[128];
			assign L0_C[130] = L0_A[0] & L0_B[130] ^ L0_A[1] & L0_B[129];
			assign L0_C[131] = L0_A[0] & L0_B[131] ^ L0_A[1] & L0_B[130];
			assign L0_C[132] = L0_A[0] & L0_B[132] ^ L0_A[1] & L0_B[131];
			assign L0_C[133] = L0_A[0] & L0_B[133] ^ L0_A[1] & L0_B[132];
			assign L0_C[134] = L0_A[0] & L0_B[134] ^ L0_A[1] & L0_B[133];
			assign L0_C[135] = L0_A[0] & L0_B[135] ^ L0_A[1] & L0_B[134];
			assign L0_C[136] = L0_A[0] & L0_B[136] ^ L0_A[1] & L0_B[135];
			assign L0_C[137] = L0_A[0] & L0_B[137] ^ L0_A[1] & L0_B[136];
			assign L0_C[138] = L0_A[0] & L0_B[138] ^ L0_A[1] & L0_B[137];
			assign L0_C[139] = L0_A[0] & L0_B[139] ^ L0_A[1] & L0_B[138];
			assign L0_C[140] = L0_A[0] & L0_B[140] ^ L0_A[1] & L0_B[139];
			assign L0_C[141] = L0_A[0] & L0_B[141] ^ L0_A[1] & L0_B[140];
			assign L0_C[142] = L0_A[0] & L0_B[142] ^ L0_A[1] & L0_B[141];
			assign L0_C[143] = L0_A[0] & L0_B[143] ^ L0_A[1] & L0_B[142];
			assign L0_C[144] = L0_A[0] & L0_B[144] ^ L0_A[1] & L0_B[143];
			assign L0_C[145] = L0_A[0] & L0_B[145] ^ L0_A[1] & L0_B[144];
			assign L0_C[146] = L0_A[0] & L0_B[146] ^ L0_A[1] & L0_B[145];
			assign L0_C[147] = L0_A[0] & L0_B[147] ^ L0_A[1] & L0_B[146];
			assign L0_C[148] = L0_A[0] & L0_B[148] ^ L0_A[1] & L0_B[147];
			assign L0_C[149] = L0_A[0] & L0_B[149] ^ L0_A[1] & L0_B[148];
			assign L0_C[150] = L0_A[0] & L0_B[150] ^ L0_A[1] & L0_B[149];
			assign L0_C[151] = L0_A[0] & L0_B[151] ^ L0_A[1] & L0_B[150];
			assign L0_C[152] = L0_A[0] & L0_B[152] ^ L0_A[1] & L0_B[151];
			assign L0_C[153] = L0_A[0] & L0_B[153] ^ L0_A[1] & L0_B[152];
			assign L0_C[154] = L0_A[0] & L0_B[154] ^ L0_A[1] & L0_B[153];
			assign L0_C[155] = L0_A[0] & L0_B[155] ^ L0_A[1] & L0_B[154];
			assign L0_C[156] = L0_A[0] & L0_B[156] ^ L0_A[1] & L0_B[155];
			assign L0_C[157] = L0_A[0] & L0_B[157] ^ L0_A[1] & L0_B[156];
			assign L0_C[158] = L0_A[0] & L0_B[158] ^ L0_A[1] & L0_B[157];
			assign L0_C[159] = L0_A[0] & L0_B[159] ^ L0_A[1] & L0_B[158];
			assign L0_C[160] = L0_A[0] & L0_B[160] ^ L0_A[1] & L0_B[159];
			assign L0_C[161] = L0_A[0] & L0_B[161] ^ L0_A[1] & L0_B[160];
			assign L0_C[162] = L0_A[0] & L0_B[162] ^ L0_A[1] & L0_B[161];
			assign L0_C[163] = L0_A[1] & L0_B[162];
			
		endmodule
