//reduRED245_c[tion 245bits
//April 21, 2009
//Yu Zhang
//yu.zhang100@gmail.com
//verified: y
													module reduction245(RED245_c, RED245_r);  
  														 input   [244:0]RED245_c;
  														 output  [162:0]RED245_r;
 								 
 								 assign RED245_r[0] = RED245_c[163]^RED245_c[0];
                 assign RED245_r[1] = RED245_c[164]^RED245_c[1];
                 assign RED245_r[2] = RED245_c[165]^RED245_c[2];
            assign RED245_r[3] = RED245_c[166]^RED245_c[3]^RED245_c[163];
            assign RED245_r[4] = RED245_c[167]^RED245_c[4]^RED245_c[164];
            assign RED245_r[5] = RED245_c[168]^RED245_c[5]^RED245_c[165];
       	assign RED245_r[6] = RED245_c[169]^RED245_c[6]^RED245_c[166]^RED245_c[163];
  			assign RED245_r[7] = RED245_c[170]^RED245_c[7]^RED245_c[167]^RED245_c[164]^RED245_c[163];
  			assign RED245_r[8] = RED245_c[171]^RED245_c[8]^RED245_c[168]^RED245_c[165]^RED245_c[164];
  			assign RED245_r[9] = RED245_c[172]^RED245_c[9]^RED245_c[169]^RED245_c[166]^RED245_c[165];
 				assign RED245_r[10] = RED245_c[173]^RED245_c[10]^RED245_c[170]^RED245_c[167]^RED245_c[166];
 				assign RED245_r[11] = RED245_c[174]^RED245_c[11]^RED245_c[171]^RED245_c[168]^RED245_c[167];
        assign RED245_r[12] = RED245_c[175]^RED245_c[12]^RED245_c[172]^RED245_c[169]^RED245_c[168];
        assign RED245_r[13] = RED245_c[176]^RED245_c[13]^RED245_c[173]^RED245_c[170]^RED245_c[169];
        assign RED245_r[14] = RED245_c[177]^RED245_c[14]^RED245_c[174]^RED245_c[171]^RED245_c[170];
        assign RED245_r[15] = RED245_c[178]^RED245_c[15]^RED245_c[175]^RED245_c[172]^RED245_c[171];
        assign RED245_r[16] = RED245_c[179]^RED245_c[16]^RED245_c[176]^RED245_c[173]^RED245_c[172];
        assign RED245_r[17] = RED245_c[180]^RED245_c[17]^RED245_c[177]^RED245_c[174]^RED245_c[173];
        assign RED245_r[18] = RED245_c[181]^RED245_c[18]^RED245_c[178]^RED245_c[175]^RED245_c[174];
        assign RED245_r[19] = RED245_c[182]^RED245_c[19]^RED245_c[179]^RED245_c[176]^RED245_c[175];
        assign RED245_r[20] = RED245_c[183]^RED245_c[20]^RED245_c[180]^RED245_c[177]^RED245_c[176];
        assign RED245_r[21] = RED245_c[184]^RED245_c[21]^RED245_c[181]^RED245_c[178]^RED245_c[177];
        assign RED245_r[22] = RED245_c[185]^RED245_c[22]^RED245_c[182]^RED245_c[179]^RED245_c[178];
        assign RED245_r[23] = RED245_c[186]^RED245_c[23]^RED245_c[183]^RED245_c[180]^RED245_c[179];
        assign RED245_r[24] = RED245_c[187]^RED245_c[24]^RED245_c[184]^RED245_c[181]^RED245_c[180];
        assign RED245_r[25] = RED245_c[188]^RED245_c[25]^RED245_c[185]^RED245_c[182]^RED245_c[181];
        assign RED245_r[26] = RED245_c[189]^RED245_c[26]^RED245_c[186]^RED245_c[183]^RED245_c[182];
        assign RED245_r[27] = RED245_c[190]^RED245_c[27]^RED245_c[187]^RED245_c[184]^RED245_c[183];
        assign RED245_r[28] = RED245_c[191]^RED245_c[28]^RED245_c[188]^RED245_c[185]^RED245_c[184];
        assign RED245_r[29] = RED245_c[192]^RED245_c[29]^RED245_c[189]^RED245_c[186]^RED245_c[185];
        assign RED245_r[30] = RED245_c[193]^RED245_c[30]^RED245_c[190]^RED245_c[187]^RED245_c[186];
        assign RED245_r[31] = RED245_c[194]^RED245_c[31]^RED245_c[191]^RED245_c[188]^RED245_c[187];
        assign RED245_r[32] = RED245_c[195]^RED245_c[32]^RED245_c[192]^RED245_c[189]^RED245_c[188];
        assign RED245_r[33] = RED245_c[196]^RED245_c[33]^RED245_c[193]^RED245_c[190]^RED245_c[189];
        assign RED245_r[34] = RED245_c[197]^RED245_c[34]^RED245_c[194]^RED245_c[191]^RED245_c[190];
        assign RED245_r[35] = RED245_c[198]^RED245_c[35]^RED245_c[195]^RED245_c[192]^RED245_c[191];
        assign RED245_r[36] = RED245_c[199]^RED245_c[36]^RED245_c[196]^RED245_c[193]^RED245_c[192];
        assign RED245_r[37] = RED245_c[200]^RED245_c[37]^RED245_c[197]^RED245_c[194]^RED245_c[193];
        assign RED245_r[38] = RED245_c[201]^RED245_c[38]^RED245_c[198]^RED245_c[195]^RED245_c[194];
        assign RED245_r[39] = RED245_c[202]^RED245_c[39]^RED245_c[199]^RED245_c[196]^RED245_c[195];
        assign RED245_r[40] = RED245_c[203]^RED245_c[40]^RED245_c[200]^RED245_c[197]^RED245_c[196];
        assign RED245_r[41] = RED245_c[204]^RED245_c[41]^RED245_c[201]^RED245_c[198]^RED245_c[197];
        assign RED245_r[42] = RED245_c[205]^RED245_c[42]^RED245_c[202]^RED245_c[199]^RED245_c[198];
        assign RED245_r[43] = RED245_c[206]^RED245_c[43]^RED245_c[203]^RED245_c[200]^RED245_c[199];
        assign RED245_r[44] = RED245_c[207]^RED245_c[44]^RED245_c[204]^RED245_c[201]^RED245_c[200];
        assign RED245_r[45] = RED245_c[208]^RED245_c[45]^RED245_c[205]^RED245_c[202]^RED245_c[201];
        assign RED245_r[46] = RED245_c[209]^RED245_c[46]^RED245_c[206]^RED245_c[203]^RED245_c[202];
        assign RED245_r[47] = RED245_c[210]^RED245_c[47]^RED245_c[207]^RED245_c[204]^RED245_c[203];
        assign RED245_r[48] = RED245_c[211]^RED245_c[48]^RED245_c[208]^RED245_c[205]^RED245_c[204];
        assign RED245_r[49] = RED245_c[212]^RED245_c[49]^RED245_c[209]^RED245_c[206]^RED245_c[205];
        assign RED245_r[50] = RED245_c[213]^RED245_c[50]^RED245_c[210]^RED245_c[207]^RED245_c[206];
        assign RED245_r[51] = RED245_c[214]^RED245_c[51]^RED245_c[211]^RED245_c[208]^RED245_c[207];
        assign RED245_r[52] = RED245_c[215]^RED245_c[52]^RED245_c[212]^RED245_c[209]^RED245_c[208];
        assign RED245_r[53] = RED245_c[216]^RED245_c[53]^RED245_c[213]^RED245_c[210]^RED245_c[209];
        assign RED245_r[54] = RED245_c[217]^RED245_c[54]^RED245_c[214]^RED245_c[211]^RED245_c[210];
        assign RED245_r[55] = RED245_c[218]^RED245_c[55]^RED245_c[215]^RED245_c[212]^RED245_c[211];
        assign RED245_r[56] = RED245_c[219]^RED245_c[56]^RED245_c[216]^RED245_c[213]^RED245_c[212];
        assign RED245_r[57] = RED245_c[220]^RED245_c[57]^RED245_c[217]^RED245_c[214]^RED245_c[213];
        assign RED245_r[58] = RED245_c[221]^RED245_c[58]^RED245_c[218]^RED245_c[215]^RED245_c[214];
        assign RED245_r[59] = RED245_c[222]^RED245_c[59]^RED245_c[219]^RED245_c[216]^RED245_c[215];
        assign RED245_r[60] = RED245_c[223]^RED245_c[60]^RED245_c[220]^RED245_c[217]^RED245_c[216];
        assign RED245_r[61] = RED245_c[224]^RED245_c[61]^RED245_c[221]^RED245_c[218]^RED245_c[217];
        assign RED245_r[62] = RED245_c[225]^RED245_c[62]^RED245_c[222]^RED245_c[219]^RED245_c[218];
        assign RED245_r[63] = RED245_c[226]^RED245_c[63]^RED245_c[223]^RED245_c[220]^RED245_c[219];
        assign RED245_r[64] = RED245_c[227]^RED245_c[64]^RED245_c[224]^RED245_c[221]^RED245_c[220];
        assign RED245_r[65] = RED245_c[228]^RED245_c[65]^RED245_c[225]^RED245_c[222]^RED245_c[221];
        assign RED245_r[66] = RED245_c[229]^RED245_c[66]^RED245_c[226]^RED245_c[223]^RED245_c[222];
        assign RED245_r[67] = RED245_c[230]^RED245_c[67]^RED245_c[227]^RED245_c[224]^RED245_c[223];
        assign RED245_r[68] = RED245_c[231]^RED245_c[68]^RED245_c[228]^RED245_c[225]^RED245_c[224];
        assign RED245_r[69] = RED245_c[232]^RED245_c[69]^RED245_c[229]^RED245_c[226]^RED245_c[225];
        assign RED245_r[70] = RED245_c[233]^RED245_c[70]^RED245_c[230]^RED245_c[227]^RED245_c[226];
        assign RED245_r[71] = RED245_c[234]^RED245_c[71]^RED245_c[231]^RED245_c[228]^RED245_c[227];
        assign RED245_r[72] = RED245_c[235]^RED245_c[72]^RED245_c[232]^RED245_c[229]^RED245_c[228];
        assign RED245_r[73] = RED245_c[236]^RED245_c[73]^RED245_c[233]^RED245_c[230]^RED245_c[229];
        assign RED245_r[74] = RED245_c[237]^RED245_c[74]^RED245_c[234]^RED245_c[231]^RED245_c[230];
        assign RED245_r[75] = RED245_c[238]^RED245_c[75]^RED245_c[235]^RED245_c[232]^RED245_c[231];
        assign RED245_r[76] = RED245_c[239]^RED245_c[76]^RED245_c[236]^RED245_c[233]^RED245_c[232];
        assign RED245_r[77] = RED245_c[240]^RED245_c[77]^RED245_c[237]^RED245_c[234]^RED245_c[233];
        assign RED245_r[78] = RED245_c[241]^RED245_c[78]^RED245_c[238]^RED245_c[235]^RED245_c[234];
        assign RED245_r[79] = RED245_c[242]^RED245_c[79]^RED245_c[239]^RED245_c[236]^RED245_c[235];
        assign RED245_r[80] = RED245_c[243]^RED245_c[80]^RED245_c[240]^RED245_c[237]^RED245_c[236];
        assign RED245_r[81] = RED245_c[244]^RED245_c[81]^RED245_c[241]^RED245_c[238]^RED245_c[237];
        assign RED245_r[82] = RED245_c[82]^RED245_c[242]^RED245_c[239]^RED245_c[238];
        assign RED245_r[83] = RED245_c[83]^RED245_c[243]^RED245_c[240]^RED245_c[239];
        assign RED245_r[84] = RED245_c[84]^RED245_c[244]^RED245_c[241]^RED245_c[240];
           assign RED245_r[85] = RED245_c[85]^RED245_c[242]^RED245_c[241];
           assign RED245_r[86] = RED245_c[86]^RED245_c[243]^RED245_c[242];
           assign RED245_r[87] = RED245_c[87]^RED245_c[244]^RED245_c[243];
                assign RED245_r[88] = RED245_c[88]^RED245_c[244];
                     assign RED245_r[89] = RED245_c[89];
                     assign RED245_r[90] = RED245_c[90];
                     assign RED245_r[91] = RED245_c[91];
                     assign RED245_r[92] = RED245_c[92];
                     assign RED245_r[93] = RED245_c[93];
                     assign RED245_r[94] = RED245_c[94];
                     assign RED245_r[95] = RED245_c[95];
                     assign RED245_r[96] = RED245_c[96];
                     assign RED245_r[97] = RED245_c[97];
                     assign RED245_r[98] = RED245_c[98];
                     assign RED245_r[99] = RED245_c[99];
                    assign RED245_r[100] = RED245_c[100];
                    assign RED245_r[101] = RED245_c[101];
                    assign RED245_r[102] = RED245_c[102];
                    assign RED245_r[103] = RED245_c[103];
                    assign RED245_r[104] = RED245_c[104];
                    assign RED245_r[105] = RED245_c[105];
                    assign RED245_r[106] = RED245_c[106];
                    assign RED245_r[107] = RED245_c[107];
                    assign RED245_r[108] = RED245_c[108];
                    assign RED245_r[109] = RED245_c[109];
                    assign RED245_r[110] = RED245_c[110];
                    assign RED245_r[111] = RED245_c[111];
                    assign RED245_r[112] = RED245_c[112];
                    assign RED245_r[113] = RED245_c[113];
                    assign RED245_r[114] = RED245_c[114];
                    assign RED245_r[115] = RED245_c[115];
                    assign RED245_r[116] = RED245_c[116];
                    assign RED245_r[117] = RED245_c[117];
                    assign RED245_r[118] = RED245_c[118];
                    assign RED245_r[119] = RED245_c[119];
                    assign RED245_r[120] = RED245_c[120];
                    assign RED245_r[121] = RED245_c[121];
                    assign RED245_r[122] = RED245_c[122];
                    assign RED245_r[123] = RED245_c[123];
                    assign RED245_r[124] = RED245_c[124];
                    assign RED245_r[125] = RED245_c[125];
                    assign RED245_r[126] = RED245_c[126];
                    assign RED245_r[127] = RED245_c[127];
                    assign RED245_r[128] = RED245_c[128];
                    assign RED245_r[129] = RED245_c[129];
                    assign RED245_r[130] = RED245_c[130];
                    assign RED245_r[131] = RED245_c[131];
                    assign RED245_r[132] = RED245_c[132];
                    assign RED245_r[133] = RED245_c[133];
                    assign RED245_r[134] = RED245_c[134];
                    assign RED245_r[135] = RED245_c[135];
                    assign RED245_r[136] = RED245_c[136];
                    assign RED245_r[137] = RED245_c[137];
                    assign RED245_r[138] = RED245_c[138];
                    assign RED245_r[139] = RED245_c[139];
                    assign RED245_r[140] = RED245_c[140];
                    assign RED245_r[141] = RED245_c[141];
                    assign RED245_r[142] = RED245_c[142];
                    assign RED245_r[143] = RED245_c[143];
                    assign RED245_r[144] = RED245_c[144];
                    assign RED245_r[145] = RED245_c[145];
                    assign RED245_r[146] = RED245_c[146];
                    assign RED245_r[147] = RED245_c[147];
                    assign RED245_r[148] = RED245_c[148];
                    assign RED245_r[149] = RED245_c[149];
                    assign RED245_r[150] = RED245_c[150];
                    assign RED245_r[151] = RED245_c[151];
                    assign RED245_r[152] = RED245_c[152];
                    assign RED245_r[153] = RED245_c[153];
                    assign RED245_r[154] = RED245_c[154];
                    assign RED245_r[155] = RED245_c[155];
                    assign RED245_r[156] = RED245_c[156];
                    assign RED245_r[157] = RED245_c[157];
                    assign RED245_r[158] = RED245_c[158];
                    assign RED245_r[159] = RED245_c[159];
                    assign RED245_r[160] = RED245_c[160];
                    assign RED245_r[161] = RED245_c[161];
                    assign RED245_r[162] = RED245_c[162];
               
                endmodule
