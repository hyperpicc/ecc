//Multiplication level3 special 
//April 21, 2009
//Yu Zhang
//yu.zhang100@gmail.com
//verified: y
module level3_special(L3S_A, L3S_B, L3S_a40, L3S_C);
			input 	[169:0]L3S_A;
			input 	[162:0]L3S_B;
			input   			 L3S_a40;
			output 	[170:0]L3S_C;
			
					assign L3S_C[0] = L3S_A[0];
					assign L3S_C[1] = L3S_A[1];
					assign L3S_C[2] = L3S_A[2];
					assign L3S_C[3] = L3S_A[3];
					assign L3S_C[4] = L3S_A[4];
					assign L3S_C[5] = L3S_A[5];
					assign L3S_C[6] = L3S_A[6];
					assign L3S_C[7] = L3S_A[7];
					assign L3S_C[8] = L3S_A[8] ^ L3S_B[0] & L3S_a40;
					assign L3S_C[9] = L3S_A[9] ^ L3S_B[1] & L3S_a40;
					assign L3S_C[10] = L3S_A[10] ^ L3S_B[2] & L3S_a40;
					assign L3S_C[11] = L3S_A[11] ^ L3S_B[3] & L3S_a40;
					assign L3S_C[12] = L3S_A[12] ^ L3S_B[4] & L3S_a40;
					assign L3S_C[13] = L3S_A[13] ^ L3S_B[5] & L3S_a40;
					assign L3S_C[14] = L3S_A[14] ^ L3S_B[6] & L3S_a40;
					assign L3S_C[15] = L3S_A[15] ^ L3S_B[7] & L3S_a40;
					assign L3S_C[16] = L3S_A[16] ^ L3S_B[8] & L3S_a40;
					assign L3S_C[17] = L3S_A[17] ^ L3S_B[9] & L3S_a40;
					assign L3S_C[18] = L3S_A[18] ^ L3S_B[10] & L3S_a40;
					assign L3S_C[19] = L3S_A[19] ^ L3S_B[11] & L3S_a40;
					assign L3S_C[20] = L3S_A[20] ^ L3S_B[12] & L3S_a40;
					assign L3S_C[21] = L3S_A[21] ^ L3S_B[13] & L3S_a40;
					assign L3S_C[22] = L3S_A[22] ^ L3S_B[14] & L3S_a40;
					assign L3S_C[23] = L3S_A[23] ^ L3S_B[15] & L3S_a40;
					assign L3S_C[24] = L3S_A[24] ^ L3S_B[16] & L3S_a40;
					assign L3S_C[25] = L3S_A[25] ^ L3S_B[17] & L3S_a40;
					assign L3S_C[26] = L3S_A[26] ^ L3S_B[18] & L3S_a40;
					assign L3S_C[27] = L3S_A[27] ^ L3S_B[19] & L3S_a40;
					assign L3S_C[28] = L3S_A[28] ^ L3S_B[20] & L3S_a40;
					assign L3S_C[29] = L3S_A[29] ^ L3S_B[21] & L3S_a40;
					assign L3S_C[30] = L3S_A[30] ^ L3S_B[22] & L3S_a40;
					assign L3S_C[31] = L3S_A[31] ^ L3S_B[23] & L3S_a40;
					assign L3S_C[32] = L3S_A[32] ^ L3S_B[24] & L3S_a40;
					assign L3S_C[33] = L3S_A[33] ^ L3S_B[25] & L3S_a40;
					assign L3S_C[34] = L3S_A[34] ^ L3S_B[26] & L3S_a40;
					assign L3S_C[35] = L3S_A[35] ^ L3S_B[27] & L3S_a40;
					assign L3S_C[36] = L3S_A[36] ^ L3S_B[28] & L3S_a40;
					assign L3S_C[37] = L3S_A[37] ^ L3S_B[29] & L3S_a40;
					assign L3S_C[38] = L3S_A[38] ^ L3S_B[30] & L3S_a40;
					assign L3S_C[39] = L3S_A[39] ^ L3S_B[31] & L3S_a40;
					assign L3S_C[40] = L3S_A[40] ^ L3S_B[32] & L3S_a40;
					assign L3S_C[41] = L3S_A[41] ^ L3S_B[33] & L3S_a40;
					assign L3S_C[42] = L3S_A[42] ^ L3S_B[34] & L3S_a40;
					assign L3S_C[43] = L3S_A[43] ^ L3S_B[35] & L3S_a40;
					assign L3S_C[44] = L3S_A[44] ^ L3S_B[36] & L3S_a40;
					assign L3S_C[45] = L3S_A[45] ^ L3S_B[37] & L3S_a40;
					assign L3S_C[46] = L3S_A[46] ^ L3S_B[38] & L3S_a40;
					assign L3S_C[47] = L3S_A[47] ^ L3S_B[39] & L3S_a40;
					assign L3S_C[48] = L3S_A[48] ^ L3S_B[40] & L3S_a40;
					assign L3S_C[49] = L3S_A[49] ^ L3S_B[41] & L3S_a40;
					assign L3S_C[50] = L3S_A[50] ^ L3S_B[42] & L3S_a40;
					assign L3S_C[51] = L3S_A[51] ^ L3S_B[43] & L3S_a40;
					assign L3S_C[52] = L3S_A[52] ^ L3S_B[44] & L3S_a40;
					assign L3S_C[53] = L3S_A[53] ^ L3S_B[45] & L3S_a40;
					assign L3S_C[54] = L3S_A[54] ^ L3S_B[46] & L3S_a40;
					assign L3S_C[55] = L3S_A[55] ^ L3S_B[47] & L3S_a40;
					assign L3S_C[56] = L3S_A[56] ^ L3S_B[48] & L3S_a40;
					assign L3S_C[57] = L3S_A[57] ^ L3S_B[49] & L3S_a40;
					assign L3S_C[58] = L3S_A[58] ^ L3S_B[50] & L3S_a40;
					assign L3S_C[59] = L3S_A[59] ^ L3S_B[51] & L3S_a40;
					assign L3S_C[60] = L3S_A[60] ^ L3S_B[52] & L3S_a40;
					assign L3S_C[61] = L3S_A[61] ^ L3S_B[53] & L3S_a40;
					assign L3S_C[62] = L3S_A[62] ^ L3S_B[54] & L3S_a40;
					assign L3S_C[63] = L3S_A[63] ^ L3S_B[55] & L3S_a40;
					assign L3S_C[64] = L3S_A[64] ^ L3S_B[56] & L3S_a40;
					assign L3S_C[65] = L3S_A[65] ^ L3S_B[57] & L3S_a40;
					assign L3S_C[66] = L3S_A[66] ^ L3S_B[58] & L3S_a40;
					assign L3S_C[67] = L3S_A[67] ^ L3S_B[59] & L3S_a40;
					assign L3S_C[68] = L3S_A[68] ^ L3S_B[60] & L3S_a40;
					assign L3S_C[69] = L3S_A[69] ^ L3S_B[61] & L3S_a40;
					assign L3S_C[70] = L3S_A[70] ^ L3S_B[62] & L3S_a40;
					assign L3S_C[71] = L3S_A[71] ^ L3S_B[63] & L3S_a40;
					assign L3S_C[72] = L3S_A[72] ^ L3S_B[64] & L3S_a40;
					assign L3S_C[73] = L3S_A[73] ^ L3S_B[65] & L3S_a40;
					assign L3S_C[74] = L3S_A[74] ^ L3S_B[66] & L3S_a40;
					assign L3S_C[75] = L3S_A[75] ^ L3S_B[67] & L3S_a40;
					assign L3S_C[76] = L3S_A[76] ^ L3S_B[68] & L3S_a40;
					assign L3S_C[77] = L3S_A[77] ^ L3S_B[69] & L3S_a40;
					assign L3S_C[78] = L3S_A[78] ^ L3S_B[70] & L3S_a40;
					assign L3S_C[79] = L3S_A[79] ^ L3S_B[71] & L3S_a40;
					assign L3S_C[80] = L3S_A[80] ^ L3S_B[72] & L3S_a40;
					assign L3S_C[81] = L3S_A[81] ^ L3S_B[73] & L3S_a40;
					assign L3S_C[82] = L3S_A[82] ^ L3S_B[74] & L3S_a40;
					assign L3S_C[83] = L3S_A[83] ^ L3S_B[75] & L3S_a40;
					assign L3S_C[84] = L3S_A[84] ^ L3S_B[76] & L3S_a40;
					assign L3S_C[85] = L3S_A[85] ^ L3S_B[77] & L3S_a40;
					assign L3S_C[86] = L3S_A[86] ^ L3S_B[78] & L3S_a40;
					assign L3S_C[87] = L3S_A[87] ^ L3S_B[79] & L3S_a40;
					assign L3S_C[88] = L3S_A[88] ^ L3S_B[80] & L3S_a40;
					assign L3S_C[89] = L3S_A[89] ^ L3S_B[81] & L3S_a40;
					assign L3S_C[90] = L3S_A[90] ^ L3S_B[82] & L3S_a40;
					assign L3S_C[91] = L3S_A[91] ^ L3S_B[83] & L3S_a40;
					assign L3S_C[92] = L3S_A[92] ^ L3S_B[84] & L3S_a40;
					assign L3S_C[93] = L3S_A[93] ^ L3S_B[85] & L3S_a40;
					assign L3S_C[94] = L3S_A[94] ^ L3S_B[86] & L3S_a40;
					assign L3S_C[95] = L3S_A[95] ^ L3S_B[87] & L3S_a40;
					assign L3S_C[96] = L3S_A[96] ^ L3S_B[88] & L3S_a40;
					assign L3S_C[97] = L3S_A[97] ^ L3S_B[89] & L3S_a40;
					assign L3S_C[98] = L3S_A[98] ^ L3S_B[90] & L3S_a40;
					assign L3S_C[99] = L3S_A[99] ^ L3S_B[91] & L3S_a40;
					assign L3S_C[100] = L3S_A[100] ^ L3S_B[92] & L3S_a40;
					assign L3S_C[101] = L3S_A[101] ^ L3S_B[93] & L3S_a40;
					assign L3S_C[102] = L3S_A[102] ^ L3S_B[94] & L3S_a40;
					assign L3S_C[103] = L3S_A[103] ^ L3S_B[95] & L3S_a40;
					assign L3S_C[104] = L3S_A[104] ^ L3S_B[96] & L3S_a40;
					assign L3S_C[105] = L3S_A[105] ^ L3S_B[97] & L3S_a40;
					assign L3S_C[106] = L3S_A[106] ^ L3S_B[98] & L3S_a40;
					assign L3S_C[107] = L3S_A[107] ^ L3S_B[99] & L3S_a40;
					assign L3S_C[108] = L3S_A[108] ^ L3S_B[100] & L3S_a40;
					assign L3S_C[109] = L3S_A[109] ^ L3S_B[101] & L3S_a40;
					assign L3S_C[110] = L3S_A[110] ^ L3S_B[102] & L3S_a40;
					assign L3S_C[111] = L3S_A[111] ^ L3S_B[103] & L3S_a40;
					assign L3S_C[112] = L3S_A[112] ^ L3S_B[104] & L3S_a40;
					assign L3S_C[113] = L3S_A[113] ^ L3S_B[105] & L3S_a40;
					assign L3S_C[114] = L3S_A[114] ^ L3S_B[106] & L3S_a40;
					assign L3S_C[115] = L3S_A[115] ^ L3S_B[107] & L3S_a40;
					assign L3S_C[116] = L3S_A[116] ^ L3S_B[108] & L3S_a40;
					assign L3S_C[117] = L3S_A[117] ^ L3S_B[109] & L3S_a40;
					assign L3S_C[118] = L3S_A[118] ^ L3S_B[110] & L3S_a40;
					assign L3S_C[119] = L3S_A[119] ^ L3S_B[111] & L3S_a40;
					assign L3S_C[120] = L3S_A[120] ^ L3S_B[112] & L3S_a40;
					assign L3S_C[121] = L3S_A[121] ^ L3S_B[113] & L3S_a40;
					assign L3S_C[122] = L3S_A[122] ^ L3S_B[114] & L3S_a40;
					assign L3S_C[123] = L3S_A[123] ^ L3S_B[115] & L3S_a40;
					assign L3S_C[124] = L3S_A[124] ^ L3S_B[116] & L3S_a40;
					assign L3S_C[125] = L3S_A[125] ^ L3S_B[117] & L3S_a40;
					assign L3S_C[126] = L3S_A[126] ^ L3S_B[118] & L3S_a40;
					assign L3S_C[127] = L3S_A[127] ^ L3S_B[119] & L3S_a40;
					assign L3S_C[128] = L3S_A[128] ^ L3S_B[120] & L3S_a40;
					assign L3S_C[129] = L3S_A[129] ^ L3S_B[121] & L3S_a40;
					assign L3S_C[130] = L3S_A[130] ^ L3S_B[122] & L3S_a40;
					assign L3S_C[131] = L3S_A[131] ^ L3S_B[123] & L3S_a40;
					assign L3S_C[132] = L3S_A[132] ^ L3S_B[124] & L3S_a40;
					assign L3S_C[133] = L3S_A[133] ^ L3S_B[125] & L3S_a40;
					assign L3S_C[134] = L3S_A[134] ^ L3S_B[126] & L3S_a40;
					assign L3S_C[135] = L3S_A[135] ^ L3S_B[127] & L3S_a40;
					assign L3S_C[136] = L3S_A[136] ^ L3S_B[128] & L3S_a40;
					assign L3S_C[137] = L3S_A[137] ^ L3S_B[129] & L3S_a40;
					assign L3S_C[138] = L3S_A[138] ^ L3S_B[130] & L3S_a40;
					assign L3S_C[139] = L3S_A[139] ^ L3S_B[131] & L3S_a40;
					assign L3S_C[140] = L3S_A[140] ^ L3S_B[132] & L3S_a40;
					assign L3S_C[141] = L3S_A[141] ^ L3S_B[133] & L3S_a40;
					assign L3S_C[142] = L3S_A[142] ^ L3S_B[134] & L3S_a40;
					assign L3S_C[143] = L3S_A[143] ^ L3S_B[135] & L3S_a40;
					assign L3S_C[144] = L3S_A[144] ^ L3S_B[136] & L3S_a40;
					assign L3S_C[145] = L3S_A[145] ^ L3S_B[137] & L3S_a40;
					assign L3S_C[146] = L3S_A[146] ^ L3S_B[138] & L3S_a40;
					assign L3S_C[147] = L3S_A[147] ^ L3S_B[139] & L3S_a40;
					assign L3S_C[148] = L3S_A[148] ^ L3S_B[140] & L3S_a40;
					assign L3S_C[149] = L3S_A[149] ^ L3S_B[141] & L3S_a40;
					assign L3S_C[150] = L3S_A[150] ^ L3S_B[142] & L3S_a40;
					assign L3S_C[151] = L3S_A[151] ^ L3S_B[143] & L3S_a40;
					assign L3S_C[152] = L3S_A[152] ^ L3S_B[144] & L3S_a40;
					assign L3S_C[153] = L3S_A[153] ^ L3S_B[145] & L3S_a40;
					assign L3S_C[154] = L3S_A[154] ^ L3S_B[146] & L3S_a40;
					assign L3S_C[155] = L3S_A[155] ^ L3S_B[147] & L3S_a40;
					assign L3S_C[156] = L3S_A[156] ^ L3S_B[148] & L3S_a40;
					assign L3S_C[157] = L3S_A[157] ^ L3S_B[149] & L3S_a40;
					assign L3S_C[158] = L3S_A[158] ^ L3S_B[150] & L3S_a40;
					assign L3S_C[159] = L3S_A[159] ^ L3S_B[151] & L3S_a40;
					assign L3S_C[160] = L3S_A[160] ^ L3S_B[152] & L3S_a40;
					assign L3S_C[161] = L3S_A[161] ^ L3S_B[153] & L3S_a40;
					assign L3S_C[162] = L3S_A[162] ^ L3S_B[154] & L3S_a40;
					assign L3S_C[163] = L3S_A[163] ^ L3S_B[155] & L3S_a40;
					assign L3S_C[164] = L3S_A[164] ^ L3S_B[156] & L3S_a40;
					assign L3S_C[165] = L3S_A[165] ^ L3S_B[157] & L3S_a40;
					assign L3S_C[166] = L3S_A[166] ^ L3S_B[158] & L3S_a40;
					assign L3S_C[167] = L3S_A[167] ^ L3S_B[159] & L3S_a40;
					assign L3S_C[168] = L3S_A[168] ^ L3S_B[160] & L3S_a40;
					assign L3S_C[169] = L3S_A[169] ^ L3S_B[161] & L3S_a40;
					assign L3S_C[170] = L3S_B[162] & L3S_a40;

			
		endmodule
			
