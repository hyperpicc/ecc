//adder
//April 27, 2009
//Yu Zhang
//yu.zhang100@gmail.com

module adder(ADD_A, ADD_B, ADD_R);
input [162:0]ADD_A;
input [162:0]ADD_B;
output [162:0]ADD_R;

wire [162:0]ADD_A;
wire [162:0]ADD_B;
wire [162:0]ADD_R;

		assign ADD_R[0] = ADD_A[0] ^ ADD_B[0];
		assign ADD_R[1] = ADD_A[1] ^ ADD_B[1];
		assign ADD_R[2] = ADD_A[2] ^ ADD_B[2];
		assign ADD_R[3] = ADD_A[3] ^ ADD_B[3];
		assign ADD_R[4] = ADD_A[4] ^ ADD_B[4];
		assign ADD_R[5] = ADD_A[5] ^ ADD_B[5];
		assign ADD_R[6] = ADD_A[6] ^ ADD_B[6];
		assign ADD_R[7] = ADD_A[7] ^ ADD_B[7];
		assign ADD_R[8] = ADD_A[8] ^ ADD_B[8];
		assign ADD_R[9] = ADD_A[9] ^ ADD_B[9];
		assign ADD_R[10] = ADD_A[10] ^ ADD_B[10];
		assign ADD_R[11] = ADD_A[11] ^ ADD_B[11];
		assign ADD_R[12] = ADD_A[12] ^ ADD_B[12];
		assign ADD_R[13] = ADD_A[13] ^ ADD_B[13];
		assign ADD_R[14] = ADD_A[14] ^ ADD_B[14];
		assign ADD_R[15] = ADD_A[15] ^ ADD_B[15];
		assign ADD_R[16] = ADD_A[16] ^ ADD_B[16];
		assign ADD_R[17] = ADD_A[17] ^ ADD_B[17];
		assign ADD_R[18] = ADD_A[18] ^ ADD_B[18];
		assign ADD_R[19] = ADD_A[19] ^ ADD_B[19];
		assign ADD_R[20] = ADD_A[20] ^ ADD_B[20];
		assign ADD_R[21] = ADD_A[21] ^ ADD_B[21];
		assign ADD_R[22] = ADD_A[22] ^ ADD_B[22];
		assign ADD_R[23] = ADD_A[23] ^ ADD_B[23];
		assign ADD_R[24] = ADD_A[24] ^ ADD_B[24];
		assign ADD_R[25] = ADD_A[25] ^ ADD_B[25];
		assign ADD_R[26] = ADD_A[26] ^ ADD_B[26];
		assign ADD_R[27] = ADD_A[27] ^ ADD_B[27];
		assign ADD_R[28] = ADD_A[28] ^ ADD_B[28];
		assign ADD_R[29] = ADD_A[29] ^ ADD_B[29];
		assign ADD_R[30] = ADD_A[30] ^ ADD_B[30];
		assign ADD_R[31] = ADD_A[31] ^ ADD_B[31];
		assign ADD_R[32] = ADD_A[32] ^ ADD_B[32];
		assign ADD_R[33] = ADD_A[33] ^ ADD_B[33];
		assign ADD_R[34] = ADD_A[34] ^ ADD_B[34];
		assign ADD_R[35] = ADD_A[35] ^ ADD_B[35];
		assign ADD_R[36] = ADD_A[36] ^ ADD_B[36];
		assign ADD_R[37] = ADD_A[37] ^ ADD_B[37];
		assign ADD_R[38] = ADD_A[38] ^ ADD_B[38];
		assign ADD_R[39] = ADD_A[39] ^ ADD_B[39];
		assign ADD_R[40] = ADD_A[40] ^ ADD_B[40];
		assign ADD_R[41] = ADD_A[41] ^ ADD_B[41];
		assign ADD_R[42] = ADD_A[42] ^ ADD_B[42];
		assign ADD_R[43] = ADD_A[43] ^ ADD_B[43];
		assign ADD_R[44] = ADD_A[44] ^ ADD_B[44];
		assign ADD_R[45] = ADD_A[45] ^ ADD_B[45];
		assign ADD_R[46] = ADD_A[46] ^ ADD_B[46];
		assign ADD_R[47] = ADD_A[47] ^ ADD_B[47];
		assign ADD_R[48] = ADD_A[48] ^ ADD_B[48];
		assign ADD_R[49] = ADD_A[49] ^ ADD_B[49];
		assign ADD_R[50] = ADD_A[50] ^ ADD_B[50];
		assign ADD_R[51] = ADD_A[51] ^ ADD_B[51];
		assign ADD_R[52] = ADD_A[52] ^ ADD_B[52];
		assign ADD_R[53] = ADD_A[53] ^ ADD_B[53];
		assign ADD_R[54] = ADD_A[54] ^ ADD_B[54];
		assign ADD_R[55] = ADD_A[55] ^ ADD_B[55];
		assign ADD_R[56] = ADD_A[56] ^ ADD_B[56];
		assign ADD_R[57] = ADD_A[57] ^ ADD_B[57];
		assign ADD_R[58] = ADD_A[58] ^ ADD_B[58];
		assign ADD_R[59] = ADD_A[59] ^ ADD_B[59];
		assign ADD_R[60] = ADD_A[60] ^ ADD_B[60];
		assign ADD_R[61] = ADD_A[61] ^ ADD_B[61];
		assign ADD_R[62] = ADD_A[62] ^ ADD_B[62];
		assign ADD_R[63] = ADD_A[63] ^ ADD_B[63];
		assign ADD_R[64] = ADD_A[64] ^ ADD_B[64];
		assign ADD_R[65] = ADD_A[65] ^ ADD_B[65];
		assign ADD_R[66] = ADD_A[66] ^ ADD_B[66];
		assign ADD_R[67] = ADD_A[67] ^ ADD_B[67];
		assign ADD_R[68] = ADD_A[68] ^ ADD_B[68];
		assign ADD_R[69] = ADD_A[69] ^ ADD_B[69];
		assign ADD_R[70] = ADD_A[70] ^ ADD_B[70];
		assign ADD_R[71] = ADD_A[71] ^ ADD_B[71];
		assign ADD_R[72] = ADD_A[72] ^ ADD_B[72];
		assign ADD_R[73] = ADD_A[73] ^ ADD_B[73];
		assign ADD_R[74] = ADD_A[74] ^ ADD_B[74];
		assign ADD_R[75] = ADD_A[75] ^ ADD_B[75];
		assign ADD_R[76] = ADD_A[76] ^ ADD_B[76];
		assign ADD_R[77] = ADD_A[77] ^ ADD_B[77];
		assign ADD_R[78] = ADD_A[78] ^ ADD_B[78];
		assign ADD_R[79] = ADD_A[79] ^ ADD_B[79];
		assign ADD_R[80] = ADD_A[80] ^ ADD_B[80];
		assign ADD_R[81] = ADD_A[81] ^ ADD_B[81];
		assign ADD_R[82] = ADD_A[82] ^ ADD_B[82];
		assign ADD_R[83] = ADD_A[83] ^ ADD_B[83];
		assign ADD_R[84] = ADD_A[84] ^ ADD_B[84];
		assign ADD_R[85] = ADD_A[85] ^ ADD_B[85];
		assign ADD_R[86] = ADD_A[86] ^ ADD_B[86];
		assign ADD_R[87] = ADD_A[87] ^ ADD_B[87];
		assign ADD_R[88] = ADD_A[88] ^ ADD_B[88];
		assign ADD_R[89] = ADD_A[89] ^ ADD_B[89];
		assign ADD_R[90] = ADD_A[90] ^ ADD_B[90];
		assign ADD_R[91] = ADD_A[91] ^ ADD_B[91];
		assign ADD_R[92] = ADD_A[92] ^ ADD_B[92];
		assign ADD_R[93] = ADD_A[93] ^ ADD_B[93];
		assign ADD_R[94] = ADD_A[94] ^ ADD_B[94];
		assign ADD_R[95] = ADD_A[95] ^ ADD_B[95];
		assign ADD_R[96] = ADD_A[96] ^ ADD_B[96];
		assign ADD_R[97] = ADD_A[97] ^ ADD_B[97];
		assign ADD_R[98] = ADD_A[98] ^ ADD_B[98];
		assign ADD_R[99] = ADD_A[99] ^ ADD_B[99];
		assign ADD_R[100] = ADD_A[100] ^ ADD_B[100];
		assign ADD_R[101] = ADD_A[101] ^ ADD_B[101];
		assign ADD_R[102] = ADD_A[102] ^ ADD_B[102];
		assign ADD_R[103] = ADD_A[103] ^ ADD_B[103];
		assign ADD_R[104] = ADD_A[104] ^ ADD_B[104];
		assign ADD_R[105] = ADD_A[105] ^ ADD_B[105];
		assign ADD_R[106] = ADD_A[106] ^ ADD_B[106];
		assign ADD_R[107] = ADD_A[107] ^ ADD_B[107];
		assign ADD_R[108] = ADD_A[108] ^ ADD_B[108];
		assign ADD_R[109] = ADD_A[109] ^ ADD_B[109];
		assign ADD_R[110] = ADD_A[110] ^ ADD_B[110];
		assign ADD_R[111] = ADD_A[111] ^ ADD_B[111];
		assign ADD_R[112] = ADD_A[112] ^ ADD_B[112];
		assign ADD_R[113] = ADD_A[113] ^ ADD_B[113];
		assign ADD_R[114] = ADD_A[114] ^ ADD_B[114];
		assign ADD_R[115] = ADD_A[115] ^ ADD_B[115];
		assign ADD_R[116] = ADD_A[116] ^ ADD_B[116];
		assign ADD_R[117] = ADD_A[117] ^ ADD_B[117];
		assign ADD_R[118] = ADD_A[118] ^ ADD_B[118];
		assign ADD_R[119] = ADD_A[119] ^ ADD_B[119];
		assign ADD_R[120] = ADD_A[120] ^ ADD_B[120];
		assign ADD_R[121] = ADD_A[121] ^ ADD_B[121];
		assign ADD_R[122] = ADD_A[122] ^ ADD_B[122];
		assign ADD_R[123] = ADD_A[123] ^ ADD_B[123];
		assign ADD_R[124] = ADD_A[124] ^ ADD_B[124];
		assign ADD_R[125] = ADD_A[125] ^ ADD_B[125];
		assign ADD_R[126] = ADD_A[126] ^ ADD_B[126];
		assign ADD_R[127] = ADD_A[127] ^ ADD_B[127];
		assign ADD_R[128] = ADD_A[128] ^ ADD_B[128];
		assign ADD_R[129] = ADD_A[129] ^ ADD_B[129];
		assign ADD_R[130] = ADD_A[130] ^ ADD_B[130];
		assign ADD_R[131] = ADD_A[131] ^ ADD_B[131];
		assign ADD_R[132] = ADD_A[132] ^ ADD_B[132];
		assign ADD_R[133] = ADD_A[133] ^ ADD_B[133];
		assign ADD_R[134] = ADD_A[134] ^ ADD_B[134];
		assign ADD_R[135] = ADD_A[135] ^ ADD_B[135];
		assign ADD_R[136] = ADD_A[136] ^ ADD_B[136];
		assign ADD_R[137] = ADD_A[137] ^ ADD_B[137];
		assign ADD_R[138] = ADD_A[138] ^ ADD_B[138];
		assign ADD_R[139] = ADD_A[139] ^ ADD_B[139];
		assign ADD_R[140] = ADD_A[140] ^ ADD_B[140];
		assign ADD_R[141] = ADD_A[141] ^ ADD_B[141];
		assign ADD_R[142] = ADD_A[142] ^ ADD_B[142];
		assign ADD_R[143] = ADD_A[143] ^ ADD_B[143];
		assign ADD_R[144] = ADD_A[144] ^ ADD_B[144];
		assign ADD_R[145] = ADD_A[145] ^ ADD_B[145];
		assign ADD_R[146] = ADD_A[146] ^ ADD_B[146];
		assign ADD_R[147] = ADD_A[147] ^ ADD_B[147];
		assign ADD_R[148] = ADD_A[148] ^ ADD_B[148];
		assign ADD_R[149] = ADD_A[149] ^ ADD_B[149];
		assign ADD_R[150] = ADD_A[150] ^ ADD_B[150];
		assign ADD_R[151] = ADD_A[151] ^ ADD_B[151];
		assign ADD_R[152] = ADD_A[152] ^ ADD_B[152];
		assign ADD_R[153] = ADD_A[153] ^ ADD_B[153];
		assign ADD_R[154] = ADD_A[154] ^ ADD_B[154];
		assign ADD_R[155] = ADD_A[155] ^ ADD_B[155];
		assign ADD_R[156] = ADD_A[156] ^ ADD_B[156];
		assign ADD_R[157] = ADD_A[157] ^ ADD_B[157];
		assign ADD_R[158] = ADD_A[158] ^ ADD_B[158];
		assign ADD_R[159] = ADD_A[159] ^ ADD_B[159];
		assign ADD_R[160] = ADD_A[160] ^ ADD_B[160];
		assign ADD_R[161] = ADD_A[161] ^ ADD_B[161];
		assign ADD_R[162] = ADD_A[162] ^ ADD_B[162];

endmodule
