`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: U of S
// Engineer: Yu Zhang

//yu.zhang100@gmail.com
// 
// Create Date:    06:37:13 06/07/2009 
// Design Name:    ecc_yop_tb
// Module Name:     ecc_yop_tb
// Project Name:   ECC Multi-Core Porcessor
// Target Devices: V4
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
// Verfified: N
//////////////////////////////////////////////////////////////////////////////////
module ecc_tb;
reg clk;
reg rst;
reg enable;

reg [162:0]din;
wire [162:0]dx;
wire [162:0]dy;
wire done;

//reg reg_rst;
//reg reg_enable;

//reg [162:0]reg_din;

wire bingo_x;
wire bingo_y;



assign bingo_x =								(dx == {3'b  001,
											 10'b	1101110011,
											 10'b 1011101111,
											 10'b 1111000111,
											 10'b 0101110001,
											 10'b 1100111110,
											 10'b 0010100011,
											 10'b 1000011000,
											 10'b 1000110011,
											 10'b 1110001001,
											 10'b 1100111111,
											 10'b 1110001000,
											 10'b 1000111100,
											 10'b 1001110001,
											 10'b 1010100110,
											 10'b 1110011110,
											 10'b 1000000111	
											 }
									)? 1:0;
									
									
assign bingo_y = (dy == {3'b 001,
											10'b 0100101100,
											10'b 1111011100,
											10'b 0001000100,
											10'b 1101001100,
											10'b 0101101001,
											10'b 1110111011,
											10'b 0010100011,
											10'b 1111000101,
											10'b 0101101010,
											10'b 0100111110,
											10'b 1100111100,
											10'b 1110100111,
											10'b 1101011011,
											10'b 0010000101,
											10'b 0101010101,
											10'b 1001011101
											} );
								

											 
//always@(posedge clk)
//	begin
//		reg_rst <= rst;
//		reg_enable <= enable;
//
//		reg_din <= din;
//	end
	
//ecc_top ecc_top_ins(clk, reg_rst,  done,reg_enable, dx, dy, reg_din);
//ecc_top ecc_top_ins(clk, reg_rst, reg_enable, reg_din, dx, dy, done);
ecc ecc_ins(.clk(clk), .rst(rst) , .enable(enable), .din(din), .dx(dx), .dy(dy), .done(done));


always
	#2.70 clk = ~clk;
	

initial
	begin
	
   
		clk = 1'b0;
		rst = 1'b1;
		enable = 1'b0;

		din = 163'd0;
		#27.0
		
		rst = 1'b0;
		#5.4
		#5.4
		#5.4 
		#5.4 
		#5.4  
		rst = 1'b1;
		
		#27.0//x

			enable = 1'b1;
			din = { 10'b 0111111000,
							10'b 0111010111,
							10'b 0100001011,
							10'b 0001010000,
							10'b 1101010001,
							10'b 0110101010,
							10'b 1111110101,
							10'b 0000010011,
							10'b 0010001000,
							10'b 1011010001,
							10'b 1010100100,
							10'b 1100101000,
							10'b 1100011011,
							10'b 1111010000,
							10'b 0110100001,
							10'b 1111000110,
							3'b 110
			};
		
		#5.4
		enable = 1'b1;//y
		din = { 10'b 0001101010,
						10'b 1000111111,
						10'b 0111100011,
						10'b 0110001110,
						10'b 0011010000,
						10'b 0000010010,
						10'b 1001111101,
						10'b 0001011001,
						10'b 1011101010,
						10'b 1010001011,
						10'b 0110001000,
						10'b 1110001011,
						10'b 1000000110,
						10'b 0011110010,
						10'b 1110011001,
						10'b 0010011110,
						3'b 001
						};
		#5.4
		enable = 1'b1;//k
		din = {3'b101,
			   10'b 1010101010,
			   10'b 1110101010,
			   10'b 1010001010,
			   10'b 1111101011,
			   10'b 1010101011,
			   10'b 0010101010,
			   10'b 1010101000,
			   10'b 1111001000,
			   10'b 0010101001,
			   10'b 1010101010,
			   10'b 1010101110,
			   10'b 1010101111,
			   10'b 0110101010,
			   10'b 1010001110,
			   10'b 1010101011,
			   10'b 1011101011
			   };	
		
		#5.4
		enable =1'b1;//b
						din = { 10'b 0100000101,
						10'b 0011000000,
						10'b 0011001000,
						10'b 0011110111,
						10'b 0001100100,
						10'b 1010100111,
						10'b 1001010000,
						10'b 1010010000,
						10'b 0011110101,
						10'b 1000100000,
						10'b 1010001001,
						10'b 0111101111,
						10'b 0000111010,
						10'b 0010010100,
						10'b 0110010000,
						10'b 0010111111,
						3'b 101
						};
		#5.4
			enable = 1'b0;
	
			
		#9450 $stop;
	end			
	
endmodule
