//Multiplication level4
//April 21, 2009
//Yu Zhang
//yu.zhang100@gmail.com
//verified: y
module level5(L5_A, L5_B, L5_C);
			input 	[193:0]L5_A;
			input 	[170:0]L5_B;
			output 	[202:0]L5_C;
			
			assign L5_C[0] = L5_A[0];
			assign L5_C[1] = L5_A[1];
			assign L5_C[2] = L5_A[2];
			assign L5_C[3] = L5_A[3];
			assign L5_C[4] = L5_A[4];
			assign L5_C[5] = L5_A[5];
			assign L5_C[6] = L5_A[6];
			assign L5_C[7] = L5_A[7];
			assign L5_C[8] = L5_A[8];
			assign L5_C[9] = L5_A[9];
			assign L5_C[10] = L5_A[10];
			assign L5_C[11] = L5_A[11];
			assign L5_C[12] = L5_A[12];
			assign L5_C[13] = L5_A[13];
			assign L5_C[14] = L5_A[14];
			assign L5_C[15] = L5_A[15];
			assign L5_C[16] = L5_A[16];
			assign L5_C[17] = L5_A[17];
			assign L5_C[18] = L5_A[18];
			assign L5_C[19] = L5_A[19];
			assign L5_C[20] = L5_A[20];
			assign L5_C[21] = L5_A[21];
			assign L5_C[22] = L5_A[22];
			assign L5_C[23] = L5_A[23];
			assign L5_C[24] = L5_A[24];
			assign L5_C[25] = L5_A[25];
			assign L5_C[26] = L5_A[26];
			assign L5_C[27] = L5_A[27];
			assign L5_C[28] = L5_A[28];
			assign L5_C[29] = L5_A[29];
			assign L5_C[30] = L5_A[30];
			assign L5_C[31] = L5_A[31];
			
			assign L5_C[32] = L5_A[32] ^ L5_B[0];
			assign L5_C[33] = L5_A[33] ^ L5_B[1];
			assign L5_C[34] = L5_A[34] ^ L5_B[2];
			assign L5_C[35] = L5_A[35] ^ L5_B[3];
			assign L5_C[36] = L5_A[36] ^ L5_B[4];
			assign L5_C[37] = L5_A[37] ^ L5_B[5];
			assign L5_C[38] = L5_A[38] ^ L5_B[6];
			assign L5_C[39] = L5_A[39] ^ L5_B[7];
			assign L5_C[40] = L5_A[40] ^ L5_B[8];
			assign L5_C[41] = L5_A[41] ^ L5_B[9];
			assign L5_C[42] = L5_A[42] ^ L5_B[10];
			assign L5_C[43] = L5_A[43] ^ L5_B[11];
			assign L5_C[44] = L5_A[44] ^ L5_B[12];
			assign L5_C[45] = L5_A[45] ^ L5_B[13];
			assign L5_C[46] = L5_A[46] ^ L5_B[14];
			assign L5_C[47] = L5_A[47] ^ L5_B[15];
			assign L5_C[48] = L5_A[48] ^ L5_B[16];
			assign L5_C[49] = L5_A[49] ^ L5_B[17];
			assign L5_C[50] = L5_A[50] ^ L5_B[18];
			assign L5_C[51] = L5_A[51] ^ L5_B[19];
			assign L5_C[52] = L5_A[52] ^ L5_B[20];
			assign L5_C[53] = L5_A[53] ^ L5_B[21];
			assign L5_C[54] = L5_A[54] ^ L5_B[22];
			assign L5_C[55] = L5_A[55] ^ L5_B[23];
			assign L5_C[56] = L5_A[56] ^ L5_B[24];
			assign L5_C[57] = L5_A[57] ^ L5_B[25];
			assign L5_C[58] = L5_A[58] ^ L5_B[26];
			assign L5_C[59] = L5_A[59] ^ L5_B[27];
			assign L5_C[60] = L5_A[60] ^ L5_B[28];
			assign L5_C[61] = L5_A[61] ^ L5_B[29];
			assign L5_C[62] = L5_A[62] ^ L5_B[30];
			assign L5_C[63] = L5_A[63] ^ L5_B[31];
			assign L5_C[64] = L5_A[64] ^ L5_B[32];
			assign L5_C[65] = L5_A[65] ^ L5_B[33];
			assign L5_C[66] = L5_A[66] ^ L5_B[34];
			assign L5_C[67] = L5_A[67] ^ L5_B[35];
			assign L5_C[68] = L5_A[68] ^ L5_B[36];
			assign L5_C[69] = L5_A[69] ^ L5_B[37];
			assign L5_C[70] = L5_A[70] ^ L5_B[38];
			assign L5_C[71] = L5_A[71] ^ L5_B[39];
			assign L5_C[72] = L5_A[72] ^ L5_B[40];
			assign L5_C[73] = L5_A[73] ^ L5_B[41];
			assign L5_C[74] = L5_A[74] ^ L5_B[42];
			assign L5_C[75] = L5_A[75] ^ L5_B[43];
			assign L5_C[76] = L5_A[76] ^ L5_B[44];
			assign L5_C[77] = L5_A[77] ^ L5_B[45];
			assign L5_C[78] = L5_A[78] ^ L5_B[46];
			assign L5_C[79] = L5_A[79] ^ L5_B[47];
			assign L5_C[80] = L5_A[80] ^ L5_B[48];
			assign L5_C[81] = L5_A[81] ^ L5_B[49];
			assign L5_C[82] = L5_A[82] ^ L5_B[50];
			assign L5_C[83] = L5_A[83] ^ L5_B[51];
			assign L5_C[84] = L5_A[84] ^ L5_B[52];
			assign L5_C[85] = L5_A[85] ^ L5_B[53];
			assign L5_C[86] = L5_A[86] ^ L5_B[54];
			assign L5_C[87] = L5_A[87] ^ L5_B[55];
			assign L5_C[88] = L5_A[88] ^ L5_B[56];
			assign L5_C[89] = L5_A[89] ^ L5_B[57];
			assign L5_C[90] = L5_A[90] ^ L5_B[58];
			assign L5_C[91] = L5_A[91] ^ L5_B[59];
			assign L5_C[92] = L5_A[92] ^ L5_B[60];
			assign L5_C[93] = L5_A[93] ^ L5_B[61];
			assign L5_C[94] = L5_A[94] ^ L5_B[62];
			assign L5_C[95] = L5_A[95] ^ L5_B[63];
			assign L5_C[96] = L5_A[96] ^ L5_B[64];
			assign L5_C[97] = L5_A[97] ^ L5_B[65];
			assign L5_C[98] = L5_A[98] ^ L5_B[66];
			assign L5_C[99] = L5_A[99] ^ L5_B[67];
			assign L5_C[100] = L5_A[100] ^ L5_B[68];
			assign L5_C[101] = L5_A[101] ^ L5_B[69];
			assign L5_C[102] = L5_A[102] ^ L5_B[70];
			assign L5_C[103] = L5_A[103] ^ L5_B[71];
			assign L5_C[104] = L5_A[104] ^ L5_B[72];
			assign L5_C[105] = L5_A[105] ^ L5_B[73];
			assign L5_C[106] = L5_A[106] ^ L5_B[74];
			assign L5_C[107] = L5_A[107] ^ L5_B[75];
			assign L5_C[108] = L5_A[108] ^ L5_B[76];
			assign L5_C[109] = L5_A[109] ^ L5_B[77];
			assign L5_C[110] = L5_A[110] ^ L5_B[78];
			assign L5_C[111] = L5_A[111] ^ L5_B[79];
			assign L5_C[112] = L5_A[112] ^ L5_B[80];
			assign L5_C[113] = L5_A[113] ^ L5_B[81];
			assign L5_C[114] = L5_A[114] ^ L5_B[82];
			assign L5_C[115] = L5_A[115] ^ L5_B[83];
			assign L5_C[116] = L5_A[116] ^ L5_B[84];
			assign L5_C[117] = L5_A[117] ^ L5_B[85];
			assign L5_C[118] = L5_A[118] ^ L5_B[86];
			assign L5_C[119] = L5_A[119] ^ L5_B[87];
			assign L5_C[120] = L5_A[120] ^ L5_B[88];
			assign L5_C[121] = L5_A[121] ^ L5_B[89];
			assign L5_C[122] = L5_A[122] ^ L5_B[90];
			assign L5_C[123] = L5_A[123] ^ L5_B[91];
			assign L5_C[124] = L5_A[124] ^ L5_B[92];
			assign L5_C[125] = L5_A[125] ^ L5_B[93];
			assign L5_C[126] = L5_A[126] ^ L5_B[94];
			assign L5_C[127] = L5_A[127] ^ L5_B[95];
			assign L5_C[128] = L5_A[128] ^ L5_B[96];
			assign L5_C[129] = L5_A[129] ^ L5_B[97];
			assign L5_C[130] = L5_A[130] ^ L5_B[98];
			assign L5_C[131] = L5_A[131] ^ L5_B[99];
			assign L5_C[132] = L5_A[132] ^ L5_B[100];
			assign L5_C[133] = L5_A[133] ^ L5_B[101];
			assign L5_C[134] = L5_A[134] ^ L5_B[102];
			assign L5_C[135] = L5_A[135] ^ L5_B[103];
			assign L5_C[136] = L5_A[136] ^ L5_B[104];
			assign L5_C[137] = L5_A[137] ^ L5_B[105];
			assign L5_C[138] = L5_A[138] ^ L5_B[106];
			assign L5_C[139] = L5_A[139] ^ L5_B[107];
			assign L5_C[140] = L5_A[140] ^ L5_B[108];
			assign L5_C[141] = L5_A[141] ^ L5_B[109];
			assign L5_C[142] = L5_A[142] ^ L5_B[110];
			assign L5_C[143] = L5_A[143] ^ L5_B[111];
			assign L5_C[144] = L5_A[144] ^ L5_B[112];
			assign L5_C[145] = L5_A[145] ^ L5_B[113];
			assign L5_C[146] = L5_A[146] ^ L5_B[114];
			assign L5_C[147] = L5_A[147] ^ L5_B[115];
			assign L5_C[148] = L5_A[148] ^ L5_B[116];
			assign L5_C[149] = L5_A[149] ^ L5_B[117];
			assign L5_C[150] = L5_A[150] ^ L5_B[118];
			assign L5_C[151] = L5_A[151] ^ L5_B[119];
			assign L5_C[152] = L5_A[152] ^ L5_B[120];
			assign L5_C[153] = L5_A[153] ^ L5_B[121];
			assign L5_C[154] = L5_A[154] ^ L5_B[122];
			assign L5_C[155] = L5_A[155] ^ L5_B[123];
			assign L5_C[156] = L5_A[156] ^ L5_B[124];
			assign L5_C[157] = L5_A[157] ^ L5_B[125];
			assign L5_C[158] = L5_A[158] ^ L5_B[126];
			assign L5_C[159] = L5_A[159] ^ L5_B[127];
			assign L5_C[160] = L5_A[160] ^ L5_B[128];
			assign L5_C[161] = L5_A[161] ^ L5_B[129];
			assign L5_C[162] = L5_A[162] ^ L5_B[130];
			assign L5_C[163] = L5_A[163] ^ L5_B[131];
			assign L5_C[164] = L5_A[164] ^ L5_B[132];
			assign L5_C[165] = L5_A[165] ^ L5_B[133];
			assign L5_C[166] = L5_A[166] ^ L5_B[134];
			assign L5_C[167] = L5_A[167] ^ L5_B[135];
			assign L5_C[168] = L5_A[168] ^ L5_B[136];
			assign L5_C[169] = L5_A[169] ^ L5_B[137];
			assign L5_C[170] = L5_A[170] ^ L5_B[138];
			assign L5_C[171] = L5_A[171] ^ L5_B[139];
			assign L5_C[172] = L5_A[172] ^ L5_B[140];
			assign L5_C[173] = L5_A[173] ^ L5_B[141];
			assign L5_C[174] = L5_A[174] ^ L5_B[142];
			assign L5_C[175] = L5_A[175] ^ L5_B[143];
			assign L5_C[176] = L5_A[176] ^ L5_B[144];
			assign L5_C[177] = L5_A[177] ^ L5_B[145];
			assign L5_C[178] = L5_A[178] ^ L5_B[146];
			assign L5_C[179] = L5_A[179] ^ L5_B[147];
			assign L5_C[180] = L5_A[180] ^ L5_B[148];
			assign L5_C[181] = L5_A[181] ^ L5_B[149];
			assign L5_C[182] = L5_A[182] ^ L5_B[150];
			assign L5_C[183] = L5_A[183] ^ L5_B[151];
			assign L5_C[184] = L5_A[184] ^ L5_B[152];
			assign L5_C[185] = L5_A[185] ^ L5_B[153];
			assign L5_C[186] = L5_A[186] ^ L5_B[154];
			assign L5_C[187] = L5_A[187] ^ L5_B[155];
			assign L5_C[188] = L5_A[188] ^ L5_B[156];
			assign L5_C[189] = L5_A[189] ^ L5_B[157];
			assign L5_C[190] = L5_A[190] ^ L5_B[158];
			assign L5_C[191] = L5_A[191] ^ L5_B[159];
			assign L5_C[192] = L5_A[192] ^ L5_B[160];
			assign L5_C[193] = L5_A[193] ^ L5_B[161];
			assign L5_C[194] = L5_B[162];
			assign L5_C[195] = L5_B[163];
			assign L5_C[196] = L5_B[164];
			assign L5_C[197] = L5_B[165];
			assign L5_C[198] = L5_B[166];
			assign L5_C[199] = L5_B[167];
			assign L5_C[200] = L5_B[168];
			assign L5_C[201] = L5_B[169];
			assign L5_C[202] = L5_B[170];

			
		endmodule
