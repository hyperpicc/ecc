//yu.zhang100@gmail.com
module rom1(ins_addr, ins_read);
input [7:0]ins_addr;
output [20:0]ins_read;
reg [20:0]ins_read;

always@(ins_addr)
	case(ins_addr)

				8'd0 :	ins_read = 21'b000_00_00000000_00000000;
				8'd1 :	ins_read = 21'b100_10_00000011_00000010;
				8'd2 :	ins_read = 21'b000_00_00000000_00000000;
				8'd3 :	ins_read = 21'b100_01_00000011_00000010;
				8'd4 :	ins_read = 21'b010_00_10100001_00000111;//LOOP
				8'd5 :	ins_read = 21'b111_11_00000101_00000110;
				8'd6 :	ins_read = 21'b000_00_00000000_00000000;
				8'd7 :	ins_read = 21'b000_00_00000000_00000000;
				8'd8 :	ins_read = 21'b101_01_00010000_00001000;
				8'd9 :	ins_read = 21'b111_00_00000001_00000000;
				8'd10 :	ins_read = 21'b000_00_00000000_00000000;
				8'd11 :	ins_read = 21'b000_00_00000000_00000000;
				8'd12 :	ins_read = 21'b100_10_00010000_00001000;
				8'd13 :	ins_read = 21'b110_11_01000000_00000110;
				8'd14 :	ins_read = 21'b000_00_00000000_00000000;
				8'd15 :	ins_read = 21'b000_00_00000000_00000000;
				8'd16 :	ins_read = 21'b101_01_00010000_00001000;
				8'd17 :	ins_read = 21'b111_00_00000001_00000000;
				8'd18 :	ins_read = 21'b000_00_00000000_00000000;
				8'd19 :	ins_read = 21'b000_00_00000000_00000000;
				8'd20 :	ins_read = 21'b100_10_00010000_00001000;
				8'd21 :	ins_read = 21'b101_00_00000111_00000010;
				8'd22 :	ins_read = 21'b111_11_01000000_00000111;
				8'd23 :	ins_read = 21'b000_00_00000000_00000000;
				8'd24 :	ins_read = 21'b000_00_00000000_00000000;
				8'd25 :	ins_read = 21'b101_00_00010000_00000010;
				8'd26 :	ins_read = 21'b111_00_01000000_00000111;
				8'd27 :	ins_read = 21'b000_00_00000000_00000000;
				8'd28 :	ins_read = 21'b000_00_00000000_00000000;
				8'd29 :	ins_read = 21'b011_00_00000000_00010000;
				8'd30 :	ins_read = 21'b111_11_00100000_00000001;
				8'd31 :	ins_read = 21'b000_00_00000000_00000000;
				8'd32 :	ins_read = 21'b000_00_00000000_00000000;
				8'd33 :	ins_read = 21'b011_00_00000000_00010000;
				8'd34 :	ins_read = 21'b011_00_00000000_00100000;
				8'd35 :	ins_read = 21'b101_00_00000010_00100000;
				8'd36 :	ins_read = 21'b111_11_01000000_00000001;
				8'd37 :	ins_read = 21'b000_00_00000000_00000000;
				8'd38 :	ins_read = 21'b010_00_00000100_00000000;//LOOP
				8'd39 :	ins_read = 21'b011_00_00000000_00010000;
				8'd40 :	ins_read = 21'b011_00_00000000_00100000;
				8'd41 :	ins_read = 21'b111_11_00100000_00000001;
				8'd42 :	ins_read = 21'b000_00_00000000_00000000;
				8'd43 :	ins_read = 21'b010_00_00001001_00000000;//LOOP
				8'd44 :	ins_read = 21'b011_00_00000000_00010000;
				8'd45 :	ins_read = 21'b011_00_00000000_00100000;
				8'd46 :	ins_read = 21'b111_11_00100000_00000001;
				8'd47 :	ins_read = 21'b000_00_00000000_00000000;
				8'd48 :	ins_read = 21'b000_00_00000000_00000000;
				8'd49 :	ins_read = 21'b101_00_00010000_00000010;
				8'd50 :	ins_read = 21'b111_00_01000000_00000111;
				8'd51 :	ins_read = 21'b000_00_00000000_00000000;
				8'd52 :	ins_read = 21'b010_00_00010011_00000000;//LOOP
				8'd53 :	ins_read = 21'b011_00_00000000_00010000;
				8'd54 :	ins_read = 21'b011_00_00000000_00100000;
				8'd55 :	ins_read = 21'b111_11_00100000_00000001;
				8'd56 :	ins_read = 21'b000_00_00000000_00000000;
				8'd57 :	ins_read = 21'b010_00_00100111_00000000;//LOOP		
				8'd58 :	ins_read = 21'b011_00_00000000_00010000;
				8'd59 :	ins_read = 21'b011_00_00000000_00100000;
				8'd60 :	ins_read = 21'b101_00_00100000_00000010;
				8'd61 :	ins_read = 21'b111_00_01000000_00000001;
				8'd62 :	ins_read = 21'b000_00_00000000_00000000;
				8'd63 :	ins_read = 21'b000_00_00000000_00000000;
				8'd64 :	ins_read = 21'b101_00_00010000_00000010;
				8'd65 :	ins_read = 21'b111_10_01000000_00000101;
				8'd66 :	ins_read = 21'b000_00_00000000_00000000;
				8'd67 :	ins_read = 21'b000_00_00000000_00000000;
				8'd68 :	ins_read = 21'b100_00_00010000_00000011;
				8'd69 :	ins_read = 21'b111_01_01000000_00000100;
				default: ins_read = 21'b000_00_00000000_00000000;


		endcase	
	endmodule
