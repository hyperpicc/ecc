//Multiplication level1
//April 21, 2009
//Yu Zhang
//yu.zhang100@gmail.com
//verified: y
			module level1(L1_A, L1_B, L1_C);
			input 	[163:0]L1_A;
			input 	[163:0]L1_B;
			output 	[165:0]L1_C;
			
			assign L1_C[0] = L1_A[0];
			assign L1_C[1] = L1_A[1];
			assign L1_C[2] = L1_A[2] ^ L1_B[0];
			assign L1_C[3] = L1_A[3] ^ L1_B[1];
			assign L1_C[4] = L1_A[4] ^ L1_B[2];
			assign L1_C[5] = L1_A[5] ^ L1_B[3];
			assign L1_C[6] = L1_A[6] ^ L1_B[4];
			assign L1_C[7] = L1_A[7] ^ L1_B[5];
			assign L1_C[8] = L1_A[8] ^ L1_B[6];
			assign L1_C[9] = L1_A[9] ^ L1_B[7];
			assign L1_C[10] = L1_A[10] ^ L1_B[8];
			assign L1_C[11] = L1_A[11] ^ L1_B[9];
			assign L1_C[12] = L1_A[12] ^ L1_B[10];
			assign L1_C[13] = L1_A[13] ^ L1_B[11];
			assign L1_C[14] = L1_A[14] ^ L1_B[12];
			assign L1_C[15] = L1_A[15] ^ L1_B[13];
			assign L1_C[16] = L1_A[16] ^ L1_B[14];
			assign L1_C[17] = L1_A[17] ^ L1_B[15];
			assign L1_C[18] = L1_A[18] ^ L1_B[16];
			assign L1_C[19] = L1_A[19] ^ L1_B[17];
			assign L1_C[20] = L1_A[20] ^ L1_B[18];
			assign L1_C[21] = L1_A[21] ^ L1_B[19];
			assign L1_C[22] = L1_A[22] ^ L1_B[20];
			assign L1_C[23] = L1_A[23] ^ L1_B[21];
			assign L1_C[24] = L1_A[24] ^ L1_B[22];
			assign L1_C[25] = L1_A[25] ^ L1_B[23];
			assign L1_C[26] = L1_A[26] ^ L1_B[24];
			assign L1_C[27] = L1_A[27] ^ L1_B[25];
			assign L1_C[28] = L1_A[28] ^ L1_B[26];
			assign L1_C[29] = L1_A[29] ^ L1_B[27];
			assign L1_C[30] = L1_A[30] ^ L1_B[28];
			assign L1_C[31] = L1_A[31] ^ L1_B[29];
			assign L1_C[32] = L1_A[32] ^ L1_B[30];
			assign L1_C[33] = L1_A[33] ^ L1_B[31];
			assign L1_C[34] = L1_A[34] ^ L1_B[32];
			assign L1_C[35] = L1_A[35] ^ L1_B[33];
			assign L1_C[36] = L1_A[36] ^ L1_B[34];
			assign L1_C[37] = L1_A[37] ^ L1_B[35];
			assign L1_C[38] = L1_A[38] ^ L1_B[36];
			assign L1_C[39] = L1_A[39] ^ L1_B[37];
			assign L1_C[40] = L1_A[40] ^ L1_B[38];
			assign L1_C[41] = L1_A[41] ^ L1_B[39];
			assign L1_C[42] = L1_A[42] ^ L1_B[40];
			assign L1_C[43] = L1_A[43] ^ L1_B[41];
			assign L1_C[44] = L1_A[44] ^ L1_B[42];
			assign L1_C[45] = L1_A[45] ^ L1_B[43];
			assign L1_C[46] = L1_A[46] ^ L1_B[44];
			assign L1_C[47] = L1_A[47] ^ L1_B[45];
			assign L1_C[48] = L1_A[48] ^ L1_B[46];
			assign L1_C[49] = L1_A[49] ^ L1_B[47];
			assign L1_C[50] = L1_A[50] ^ L1_B[48];
			assign L1_C[51] = L1_A[51] ^ L1_B[49];
			assign L1_C[52] = L1_A[52] ^ L1_B[50];
			assign L1_C[53] = L1_A[53] ^ L1_B[51];
			assign L1_C[54] = L1_A[54] ^ L1_B[52];
			assign L1_C[55] = L1_A[55] ^ L1_B[53];
			assign L1_C[56] = L1_A[56] ^ L1_B[54];
			assign L1_C[57] = L1_A[57] ^ L1_B[55];
			assign L1_C[58] = L1_A[58] ^ L1_B[56];
			assign L1_C[59] = L1_A[59] ^ L1_B[57];
			assign L1_C[60] = L1_A[60] ^ L1_B[58];
			assign L1_C[61] = L1_A[61] ^ L1_B[59];
			assign L1_C[62] = L1_A[62] ^ L1_B[60];
			assign L1_C[63] = L1_A[63] ^ L1_B[61];
			assign L1_C[64] = L1_A[64] ^ L1_B[62];
			assign L1_C[65] = L1_A[65] ^ L1_B[63];
			assign L1_C[66] = L1_A[66] ^ L1_B[64];
			assign L1_C[67] = L1_A[67] ^ L1_B[65];
			assign L1_C[68] = L1_A[68] ^ L1_B[66];
			assign L1_C[69] = L1_A[69] ^ L1_B[67];
			assign L1_C[70] = L1_A[70] ^ L1_B[68];
			assign L1_C[71] = L1_A[71] ^ L1_B[69];
			assign L1_C[72] = L1_A[72] ^ L1_B[70];
			assign L1_C[73] = L1_A[73] ^ L1_B[71];
			assign L1_C[74] = L1_A[74] ^ L1_B[72];
			assign L1_C[75] = L1_A[75] ^ L1_B[73];
			assign L1_C[76] = L1_A[76] ^ L1_B[74];
			assign L1_C[77] = L1_A[77] ^ L1_B[75];
			assign L1_C[78] = L1_A[78] ^ L1_B[76];
			assign L1_C[79] = L1_A[79] ^ L1_B[77];
			assign L1_C[80] = L1_A[80] ^ L1_B[78];
			assign L1_C[81] = L1_A[81] ^ L1_B[79];
			assign L1_C[82] = L1_A[82] ^ L1_B[80];
			assign L1_C[83] = L1_A[83] ^ L1_B[81];
			assign L1_C[84] = L1_A[84] ^ L1_B[82];
			assign L1_C[85] = L1_A[85] ^ L1_B[83];
			assign L1_C[86] = L1_A[86] ^ L1_B[84];
			assign L1_C[87] = L1_A[87] ^ L1_B[85];
			assign L1_C[88] = L1_A[88] ^ L1_B[86];
			assign L1_C[89] = L1_A[89] ^ L1_B[87];
			assign L1_C[90] = L1_A[90] ^ L1_B[88];
			assign L1_C[91] = L1_A[91] ^ L1_B[89];
			assign L1_C[92] = L1_A[92] ^ L1_B[90];
			assign L1_C[93] = L1_A[93] ^ L1_B[91];
			assign L1_C[94] = L1_A[94] ^ L1_B[92];
			assign L1_C[95] = L1_A[95] ^ L1_B[93];
			assign L1_C[96] = L1_A[96] ^ L1_B[94];
			assign L1_C[97] = L1_A[97] ^ L1_B[95];
			assign L1_C[98] = L1_A[98] ^ L1_B[96];
			assign L1_C[99] = L1_A[99] ^ L1_B[97];
			assign L1_C[100] = L1_A[100] ^ L1_B[98];
			assign L1_C[101] = L1_A[101] ^ L1_B[99];
			assign L1_C[102] = L1_A[102] ^ L1_B[100];
			assign L1_C[103] = L1_A[103] ^ L1_B[101];
			assign L1_C[104] = L1_A[104] ^ L1_B[102];
			assign L1_C[105] = L1_A[105] ^ L1_B[103];
			assign L1_C[106] = L1_A[106] ^ L1_B[104];
			assign L1_C[107] = L1_A[107] ^ L1_B[105];
			assign L1_C[108] = L1_A[108] ^ L1_B[106];
			assign L1_C[109] = L1_A[109] ^ L1_B[107];
			assign L1_C[110] = L1_A[110] ^ L1_B[108];
			assign L1_C[111] = L1_A[111] ^ L1_B[109];
			assign L1_C[112] = L1_A[112] ^ L1_B[110];
			assign L1_C[113] = L1_A[113] ^ L1_B[111];
			assign L1_C[114] = L1_A[114] ^ L1_B[112];
			assign L1_C[115] = L1_A[115] ^ L1_B[113];
			assign L1_C[116] = L1_A[116] ^ L1_B[114];
			assign L1_C[117] = L1_A[117] ^ L1_B[115];
			assign L1_C[118] = L1_A[118] ^ L1_B[116];
			assign L1_C[119] = L1_A[119] ^ L1_B[117];
			assign L1_C[120] = L1_A[120] ^ L1_B[118];
			assign L1_C[121] = L1_A[121] ^ L1_B[119];
			assign L1_C[122] = L1_A[122] ^ L1_B[120];
			assign L1_C[123] = L1_A[123] ^ L1_B[121];
			assign L1_C[124] = L1_A[124] ^ L1_B[122];
			assign L1_C[125] = L1_A[125] ^ L1_B[123];
			assign L1_C[126] = L1_A[126] ^ L1_B[124];
			assign L1_C[127] = L1_A[127] ^ L1_B[125];
			assign L1_C[128] = L1_A[128] ^ L1_B[126];
			assign L1_C[129] = L1_A[129] ^ L1_B[127];
			assign L1_C[130] = L1_A[130] ^ L1_B[128];
			assign L1_C[131] = L1_A[131] ^ L1_B[129];
			assign L1_C[132] = L1_A[132] ^ L1_B[130];
			assign L1_C[133] = L1_A[133] ^ L1_B[131];
			assign L1_C[134] = L1_A[134] ^ L1_B[132];
			assign L1_C[135] = L1_A[135] ^ L1_B[133];
			assign L1_C[136] = L1_A[136] ^ L1_B[134];
			assign L1_C[137] = L1_A[137] ^ L1_B[135];
			assign L1_C[138] = L1_A[138] ^ L1_B[136];
			assign L1_C[139] = L1_A[139] ^ L1_B[137];
			assign L1_C[140] = L1_A[140] ^ L1_B[138];
			assign L1_C[141] = L1_A[141] ^ L1_B[139];
			assign L1_C[142] = L1_A[142] ^ L1_B[140];
			assign L1_C[143] = L1_A[143] ^ L1_B[141];
			assign L1_C[144] = L1_A[144] ^ L1_B[142];
			assign L1_C[145] = L1_A[145] ^ L1_B[143];
			assign L1_C[146] = L1_A[146] ^ L1_B[144];
			assign L1_C[147] = L1_A[147] ^ L1_B[145];
			assign L1_C[148] = L1_A[148] ^ L1_B[146];
			assign L1_C[149] = L1_A[149] ^ L1_B[147];
			assign L1_C[150] = L1_A[150] ^ L1_B[148];
			assign L1_C[151] = L1_A[151] ^ L1_B[149];
			assign L1_C[152] = L1_A[152] ^ L1_B[150];
			assign L1_C[153] = L1_A[153] ^ L1_B[151];
			assign L1_C[154] = L1_A[154] ^ L1_B[152];
			assign L1_C[155] = L1_A[155] ^ L1_B[153];
			assign L1_C[156] = L1_A[156] ^ L1_B[154];
			assign L1_C[157] = L1_A[157] ^ L1_B[155];
			assign L1_C[158] = L1_A[158] ^ L1_B[156];
			assign L1_C[159] = L1_A[159] ^ L1_B[157];
			assign L1_C[160] = L1_A[160] ^ L1_B[158];
			assign L1_C[161] = L1_A[161] ^ L1_B[159];
			assign L1_C[162] = L1_A[162] ^ L1_B[160];
			assign L1_C[163] = L1_A[163] ^ L1_B[161];
			assign L1_C[164] = L1_B[162];
			assign L1_C[165] = L1_B[163];
		endmodule
